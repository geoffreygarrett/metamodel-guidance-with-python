�csrc.surrogate.models.ffnn
SimpleRectangularNN
q )�q}q(X   _backendqctorch.nn.backends.thnn
_get_thnn_function_backend
q)RqX   _parametersqccollections
OrderedDict
q)RqX   _buffersq	h)Rq
X   _backward_hooksqh)RqX   _forward_hooksqh)RqX   _forward_pre_hooksqh)RqX   _state_dict_hooksqh)RqX   _load_state_dict_pre_hooksqh)RqX   _modulesqh)Rq(X   fc_inqctorch.nn.modules.container
Sequential
q)�q}q(hhhh)Rqh	h)Rqhh)Rqhh)Rqhh)Rqhh)Rq hh)Rq!hh)Rq"(X   0q#ctorch.nn.modules.linear
Linear
q$)�q%}q&(hhhh)Rq'(X   weightq(ctorch._utils
_rebuild_parameter
q)ctorch._utils
_rebuild_tensor_v2
q*(ctorch.storage
_load_from_bytes
q+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889221810816qX   cpuqMnNtqQ.�]q X   94889221810816qa.n      ��h�9 �=\��<��>���v���q�>>u���60�> >�=�<���难�~ھ�~"�,<9>_�=I8���:�������j$�j2�>�Ծ;^D>��[=[�?��*�3�?T�=���>5@;�+�����>س��(<"z�>r������5�>�S��ߛ���(	?�qD>��?��W>��>�/5�C>�x�>n=>��<��H>���S�?1WV>W ��>�;��Ӿ���>�[���N�>�Q�Ѷ���Q=Q*�>���=�?�.پ艚�8z�>��x�ye=:{>������>����ݚ��?��,=j��;������=Qx�=n@>S�>g?��>��a�d =�ڽg 0>��L>�_=��K�:Kνl���:�e�>�=nnj��C��fÃ>D��>r!�>�+�����@J��_������>`�;��9>�?��vM۾j�n>5�>m��h��>WԵ>���>���>��<�y>�S	����sS�uv4��ݼ��ܾbo^>"T�=���A���ؔ>�)���� �H����>f��i5��}G�o�H=�����������<x� �u�\��yY>���*T{�
��^Ҥ���>o��>��J��@�>OK=��苾_��>�x>VD���>'�ͽmu���%>nD�=,�����~���>~)�>�?Y��>o�|>�Vn��u��R�>0�T>����h��d�ξ������?[��>�$����R=�)?|����>��>���>"���j��Dk�������6=Tʾx�=W?�ӆ�i� ����>��C�>/'ݾ4q�>C��< �����7����,�>���>` ����>�\���ُ�������>�>w��j�'��>�cؾ8ݾ4�I>�g����=�j˾ϟ�>� ����=W[�վ>��ӽ��?�Z	��>t�>����+*?�]!��>?�X�hlR�~{�=c|�=�]"����^Ҕ�j�>*-龔<�� ���[=�ξ�Mj>GZݽ:�]�W��<���=_q>�۽լ>���������f�?�s��n�>�a?II�>�iʾ�m?|%��jO>��r>�R�>I��>���S=#��>%F�<=��>�?���>�J
��8��#���>��x>"s�=��,�/-_=D;�>��>�d�>.�a5]=7��S�=>I ��P��0=m�ޝ	�EbϾ&��>����>�P�����^���&=q��_A������!��>�5?�|�=�D�VĖ>�?�>�;�>8�>@9���+>k�?��,>���>,�(��"�m��Q�JF	>۱U>� ½�ʘ��Y<<@�>�VO>��
?� ׽�@�=��]>�賾;��>��澬4���=��u��>����l>g?��V>�M�<���>6�a��ʒ�).����t_׾��s;�L>��1>F�żq,�q-Rq.K KzK�q/KK�q0�h)Rq1tq2Rq3�h)Rq4�q5Rq6X   biasq7h)h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222419936qX   cpuqKzNtqQ.�]q X   94889222419936qa.z       *%
�3H��ׁ��=;�29��UX?��¾Due=9t��隽` ?�����IϾ������澮�>Yzg�BV��x=4.�>���>�b̾��>�	�>��f ?ѳ ��9��г>���`"!?��>���h�Y�9?�=2��9�j>7�?:G���M ?��V>T~h>�y��$�>ē���xq>�֏>�ш>�?����>���>;
�>p',����>6�>ߩf>�վ����=�A_>�I�=�v�>���>��۵��!���=�>�*�>y��S>�<=�z��`�z>�6{�F�?� ��R�?��@>�gY>����Y���O�>C��ky?��>��i�i��>��>��>VSS=�)y>�A�<�	�L�v>�v>Ќ�1W?���>J�\>�g>>���]���/�>YEZ>6���V>;�f�(����.?�^�b��>
?6��>Z�>ݱ��o=�]?�?� �>�?�Ǜ=q8�q9Rq:K Kz�q;K�q<�h)Rq=tq>Rq?�h)Rq@�qARqBuh	h)RqChh)RqDhh)RqEhh)RqFhh)RqGhh)RqHhh)RqIX   trainingqJ�X   in_featuresqKKX   out_featuresqLcnumpy.core.multiarray
scalar
qMcnumpy
dtype
qNX   i8qOK K�qPRqQ(KX   <qRNNNJ����J����K tqSbCz       qT�qURqVubX   1qWctorch.nn.modules.activation
LeakyReLU
qX)�qY}qZ(hhhh)Rq[h	h)Rq\hh)Rq]hh)Rq^hh)Rq_hh)Rq`hh)Rqahh)RqbhJ�X   negative_slopeqcG?�z�G�{X   inplaceqd�ubX   2qectorch.nn.modules.dropout
Dropout
qf)�qg}qh(hhhh)Rqih	h)Rqjhh)Rqkhh)Rqlhh)Rqmhh)Rqnhh)Rqohh)RqphJ�X   pqqhMhNX   f8qrK K�qsRqt(KhRNNNJ����J����K tqubC4��H[?qv�qwRqxhd�ubX   3qyctorch.nn.modules.batchnorm
BatchNorm1d
qz)�q{}q|(hhhh)Rq}(h(h)h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222105504qX   cpuqKzNtqQ.�]q X   94889222105504qa.z       ��e?��?-}?�2p?e�?�q?a��?h��?
��?"�x?�p?T~�?���?�!v?��s?=Ǆ?�?�'w?�~y?7�?��?Yz?ds?(�x?���?oU�?C|?h�x?Z�l?"X�? �m?�?�u?�Cu?<�{?��g?��?��w?y݅?�?`�v?�ۄ?9�?J��?��j?�d�?�݂?]�{?�*s?���?�A�?�y?t��?@X~?i�?u+{?��j?kau?���?�{�?�-�?box?ĵ�?�9u?�xw?ku?^ir?�|?���?&Ɉ?�1�?U$�?(�t?p? S�?]ш?Hx�?��i?Q*�?��w?n�?��o?�3�? O�?�p?��?Aj?�O�?�Gs?0�}?dM�?�P~?	�p?�?_Om?�Pv?`��?ܳt?��b?C�s?#.�?v�y?��?~�?SDu?��?|�}?" �?k�?�w?��?*��?d�?*�?q�{?��k?3��?���?�6x?��~?��l?�{�?q~�qRq�K Kz�q�K�q��h)Rq�tq�Rq��h)Rq��q�Rq�h7h)h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222688800qX   cpuqKzNtqQ.�]q X   94889222688800qa.z       ��۽4��<��@�o
�Of�<��X=m��;�˨�많����N�<C��<�Q=r�J�m �=��0��+��^9;K����}];楽ۮ��(�<j�=�zҪ�oc׼I�ʼ�.����	��{!=vw�J�z��y��j=��=Y7c�`�=u&G<C�'=M�"=��*;��F�35��m�������7��-�{��|�<z=���=}�=��$=Ț��g :FV��r�A��8��w��<�~�<�Ц��9=�y�=�R(�¤=��=��H=�-l����<�e%��:= L=,3���=!<�=k-���S)��= hs=�qg�ZL|��1�ԑ�:l	�=mt�=���;�6e�*ǉ=�$��$��<(Uf=hR;����U�2=���֣(<�;�@�+=�' =�[�����<R��C.<j�<~����ʋ�$��;�'Լ���=�����˼|$���5��E �=Q,��@��RL8<Kh5=N=�ʍ=�r��2�;X2�q��q�Rq�K Kz�q�K�q��h)Rq�tq�Rq��h)Rq��q�Rq�uh	h)Rq�(X   running_meanq�h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889221858528qX   cpuqKzNtqQ.�]q X   94889221858528qa.z       B���ډ:u=��U�O�Ļ�>9��_P�<���>:x$>z-3>�ק���x���:���=r��> ��;%6�=��~�>��>�h�<�M3>t��>=T%:��>�ջZ�=�D?g��9?��;|�ѻ�1=WϚ=�7@;i�>�U�>��m�Yk?�=�=���=��T���u=�c���|Z<@�%>vϠ;q��=Җϻ�(>�0?��>BL"=��=���=?V?5��;+?X;��$���>��Z>��G?~J[>)�(�H;灂���-?i��>~�G�>l�>�P�~ݹ=Y𣻑��>K����?�>�Tx>c��6�|�ώ>X8Z;�dY>�@A=��.�}��>��o:�'	?x��> �>,�?�J���T'?Tj<�ꚻ��?L�)?�>
�=4+�ͱ��V>2є<5=л�3�>$�>�};�g?}:��T&j>�O�>���>�	�>V��x8�=I�?��>?K�M=�@>n@E>q��q�Rq�K Kz�q�K�q��h)Rq�tq�Rq�X   running_varq�h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222173584qX   cpuqKzNtqQ.�]q X   94889222173584qa.z       {��=Hv�=X�>���= �=*�>x �=� �=�d)>|�>ۺ>�&�=���=*��=Hn>w1>���=�>���=(�>�H>��=�>n�>���=Я0>���=(E�=��$>`��=�F>�[�=���=>>��
>m�=&Q>;�>��=�m">l>�>�=��=�>���=���=� >�4�=G>��=�L>��>�
>�>^w>f�>�a?>��=��=���=V�;>?�>�>(�>x��=���=���=$�>�>���=Oa!>��>X��=�>4��=�>���=%�	>6Y>t�>�=r��=�4>��=�$
>f5>y��=� 	>5O�=��&>�U*>�>I-#>���=iL#>ڈ�=���=��>��>�w>���=��=6��=[�>�'�=j��=��>�$>Z��=|�>@��=�>��>B%>x>���=5p>�->&1>�>�>��>q��q�Rq�K Kz�q�K�q��h)Rq�tq�Rq�X   num_batches_trackedq�h*(h+B  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
LongStorage
qX   94889222173968qX   cpuqKNtqQ.�]q X   94889222173968qa.              q��q�Rq�K ))�h)Rq�tq�Rq�uhh)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hJ�X   num_featuresq�hVX   epsq�G>�����h�X   momentumq�G?�������X   affineq��X   track_running_statsq��ubuhJ�ubX	   fc_centerq�h)�q�}q�(hhhh)Rq�h	h)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�(X   0q�h$)�q�}q�(hhhh)Rq�(h(h)h*(h+B��  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222369504qX   cpuqM$:NtqQ.�]q X   94889222369504qa.$:      �ޯ��Z��������ȼ®�=)r齡��<�w�<�1ݽ�I��ȃ����;:^m9��j�=;�O=r��:�>�<~�=9�>>�нH�~�o�4����=z�=f1�"���/廔
�=K���i�=G�=W��<.���*�6<���<��Ͻ�4]����D2�=�r���%�n��g��;�i=OE�w��=��=ڡ�:� =�N�=�d��l�v�S.��#zA=F�2���=�=CA�=��#>�<B�3�oq���M�����K����=2ƃ<
�!=j(c=��':l�>�<4#��o������q����=���=閩=��<��=;��V=��=]8Խ�t�=3#/�9
��_4�=}Ϛ=�\E<�����I:-�<�Ȣ�[��<dY��(>^V6<���<Ǆ=���X7�=[�-=.½��|�w%�R��L7>Ҫ��R��{nW��60���7=ҭ-����=�D�=9a��YQ�>lZ�� �=;�^$7=P�N=+�=R՛���+��I��q��=�c�;wO��4x����u<x��2x�<1���vU=V��=��<X������4��<w��=���>>�!���:�<Q&��)�Z8�=���;�ڽC�=�`.=�=7==�=��+=#��%��=�K|=���=���<Q��Ug=	�u=�A�=9V�Vd��W�<�n0�(諒ݿ}=6d�=�o�=����0�״ӽ�L��,�2�	U��B���J7��	�Q</�>R�N=��ܽ있=�`<:�u�������<"�>�ܑ=m�=�kཁ*��[�=kqp=���=(!�=K�=�~;�u��=��a������D=y��~��X�e=���=�r��j*=��/�Q!=<��=W8˼\��=Cn>]c�;��ҽ��ۼ�ٽD�����罕e��� G�}�8>�֔=�$����=���<9���d�=�d�=����^G���Y=�h�=���=�--��s�<4c�<����I=⊴����$����&>"W���P�J9F���D�֟����<�Q�=�.>b$q=1֯���=l9!>ɀ<�����:�<-鳼�7l�H�����л�Y�0�=�>;�e�.��=�;�d��=�,��X*˽�j���h<^�<���<2���j�=�R���u�&�;�$���9��mQ�պJ<�-ʼ�K��7�F�I,���gý�sH�p�*�o �S*��K�=}k�=�'�=�<����]n=\�<Qq�<��#�{0z�S�=���=��8�=�x�ʌv=҉������rF��:�=\C�=�h�=S��OLJ=�cj�l�����Žp�3�7�>�<�xP�<���=^Ҽ`�=z0=�r=,6�<���<��C=��T���=͔�<%<��ݽmy��H,%>�W�=kbx�,����%� ;��	�=�1=Š��_=v�b�=���=�-ŽE�p<��kx<���<<=��ѼxzK=d�/=���\=���<�hr��C���n�<ڧ����=h�=*-�=�J�=���=V�k=��Q���=�>�s<�$�Z�<��<���#w�=ܖ���4�$���/�-=<ɑ� �=��
>����*���=�&�|I�&��Y�9��+1����<�L�=Jg}�>t����=�?�=�ɻˋ>��="�'=z�лW$���fTp��'i��
:�T@��5'�%cs=�܄= �=J������\�=��%���ڽ�g�<��<���9�m=�*>4)�<l��;����r��;�=F}�=�ϗ<[��=��=�ǽ�h�;n� =�E?=�Eý$��=V�>ƥ<��<���=�G8=�����d��Uн�����=�dI�y�%=F�=����=�Ua��">!(�3�'<�ф���,�� ս{=�����ỗ�*=�+\�O�X�U��u��=�1�'(ؽ T����O<�_�=hL�=��;����<Pn��勽\��h#�=��p=���y�<���;&�#��^b=3:�R��׽�:s�H������=���=t���N�Fx�D֏=�{ҽ�kW��ͽ��=�����>������<x�%>��7=0�:6��g����=\k=��K��!>�>v�=�H߻�jf; �1=�Z�=�B�=l�>=?�F��Ȝ=�}��d;�=_��G�=��>'
�*O��I���;�G�d���۽��:�G+&=���/��8<�c=��Žn�k�����5E��,�8���*>?r�=Z_=�.Ľ54�=BKL=�Ž��=���R�'�4�&��ý�垽�����%���k�X����<��4�5{ͽe������I*�=K9��<G���i<쨞< r�<�,�=���=�y��!=S�ӽ�B׼|��<��ƾ�=��ûQJ<���U=�2:sX��1�b=�IJ�'-W=�r��a&��b>��o|Լ:�=������+�� ���=���=��=l��=�#�= ����JH=�=Q����Л=��<��<N�����>�6=>ԃ=�wY;؎���qv<hT�=��<1s���<7��M�$�<s޽S��=lZ̻aQ��f�:v\�4�*�*�1<j��<�Ͻ�>:��K��5%:��f�;+f���VϽ�� =��;��\��v������>��� �-:re�=�!�<��߽�������ݰ��������=�1��=;�;K��c��=�y��İ��n/׽Z��x|w����<�G��##j=�B�=��:5�=0��5�%�Օ���:df�=�5v�()S=�k�����=T�f<&s{�����<��<.�=��	>@��="V��<@y;Rȼ���=)���wK�==қ�ѩ�=��/��d�[=گ����N=#�����=ˢ���z����!��l=b���xA�=ԅ3���N=��>����p#<���=שb�Ż=������=�-<���e�s���8}����=ɳ/<7t߽P�j;;N���ei��Q<=�h���ߩ����=@5��+��;#k8<P�=����;��?�����
#>E,=��RN��O=/Z!<k�7��� �ei�D�˽�`��μ%�:=Ȇ�<>$'=��>vv�=��R=�2�<$�[=�c< t��{�����=�.>.�<⡯<���<f�+=�t=X�J9s4��cę:*n(>@Ub�S��Xw���af=�=��b�ΐ/=	�f=gL<bM�g� =�������<d��< sʽC�H=4} >�5w<�����ӱ����������=���<L�;'��{=��T=T
[<B1����=0:9����9;ug�=@�=�g�=|�=1��<���;"aB�����y���1�<u=>$��ɀ��-+>�`��(x=\�<���=T;������=�g���_�����;6G���B��/>�@8���?�&d�=]I����<��k=p�u=4�<�֯=��=��<-�Ѽt"����<w�h�� =�系�=���1��8>B�+��"�=�1�=��k=K�3<'#J��pi��=�j�<zG��Q�(��ȽC��� ,�=�.�=)�<`�<��9��5<#�N=H���7��=�Yར��<!�~��|M=#~�=2�<=�P�=�P�=SkY=?Y�<yL=++����=����ן=����=�e<��]<��f���;��μ
��=�03�ʒ>��n=�>ZG=�c�=~�=Ҩo=��	���ջ��s���=h*�<�<�v|����<�^�[!=v��=����U�T=�F[=�.���[���w=��=��<b�<��<�&�=�W��iL��_xB=�P�	��w�P=�V	�	0�=04�=]1����v=~�'>��k�;c�;��
�0)=g8�׬=��>Og)�䃚<ҁd=�떽�l�=x7罅��<p��W7�=���<PU2��G1�X� >���^q=G޺�5a=����Oe���X�e���uk�=D����.������)>=xO<\I����<��k�e��hN�<_� ����=�ɽ���=��I������52m<���<3���C�@=Q^z<�tM=���0@r�҆�Nm!�N[7��H���$�=ٺ�u`�:�6�u?�=�D=u�m=����R������<�> ��C >J�Ž�=��;ˬ�=S�Q��V���?�����<�o����<�z����=�Fh=��=(��=^ 7��M���u�b��2<�N�<���⫧� a��di�����M8��0�=���=���=t�;�Շ�|�<� t�-�.�/�E��=���<��=��>�������,�;��<�3�l��;�>�<0|:;�b=��>X>s�5��ͻI���:�=�h��o%��3D<��y�4;�=4Q��͢=uo�}"�=k}=N�=�5=�j�(<�����=j�>=X�Խ������x��<N��;�R�=�%����L=�q�����������>�>��=��<��Խek<?�c=zU�=5!=>NϽ���=������<7��^�=�ӽX�=N'�=]`�#B�=�<Q��=���=��=:�W=m�=��=$\��F��l���>�J����=���%ߏ�+A>�S���T�sc�N�=�_�;f�<<���x!K=���	�=�s���Ƽ�~��r�P��=��=�W	>�D<y��<oܖ�%�)�lp�<[��<���;M�_��ᘽSƼKˠ�,늼�,�=���=B�d<�B����)=61<���=��P�Q��=����
<{C=C(> ����>�>T�%=(��=ꡏ��g�=��n<��H������=�I�a[��������=�s�N�ü�m�=�%>qa��z~;�;=��轻��=G��;��;kQ`=�m��J�<R�=e��<aw�=ce���󴽿J1>��]">��=�G�ES���qȼX/>������<d�;�e ;��>��H���.���38�1Ƚ��<�=�=��!��'>�σ<n����=1�=n����ڽ#������,;H=K̢=�#F=>���'`��	:��N=/ 5��^�=�Ž��޼}#�=�Ǣ=�c��L�=���;�����s���<I����=���=��=�6���=,L�=��<����|����<�<n�_=i����o1>[��eμ-�	�A"<�"=�Z�=��y����Oc�<�
�	ؼ�p]<"=���_C���=������=��;�A=_�O����<����>�mO�������=��=PZ=9�tq5=[|Ƚ����߆��p꽜�<��U<�~7��U�=1  =P�
�5��<G�=J�=��|�=���=j��ß���R����L=��μiU�=9\�/3��*���N��p���;��<�*+=t9=Z4<mW�=�ޑ�2S�����;���=F1+=B����'ֽ��<�=N��i^�l�=�詽??������<�<��=�K}<瑧�۠=�j���<C����dw�=��/<[�I<7>=�x=/rn=�����<�*�=65�=#D�='���fj���=�ɐ:�V��>1�=��<�z�=���;A_�=ټ�=L�=n��-X=q�����6q<�j>�̸=�)ϼ!�y�_.��,ED����1n=/nj='��=Z��<��)� �>sA�=��k��=��>���<DȻx�#�����I���m׽���=�=*p߽)��8���=:~E=PG,�jo���\n�6b>�A ����<���?�t�E�p�7�=6ڋ=�������J>ل�_�<g���8�^��B����"U��a��v���=M)��Vv���·=�{<P(�=���<�='B=�K���={�h��m�=e8:=��~���Q;�v�=�h�t��\Eǽ�7�=J�<��=�9�<���)W>�s��=�v��ދ�=�5���E�=Q��< ix;!g;i3�<��=�L=
�;�=�$(=q�����=uӼ���=�>�㐽�0@=�A<��>��=Ȍ�z=>���W�s�c�<������߽�v�=u��=ލ9=~1=�>?R��<�cI�����ɭ�=*�黰��҆�=~p�=�?�<:I�?_~��&�;�nսy�Y=��f��L�=G )=�=��"=�0�%��<Z�k����=8��=����#��^T��e�<_�<�WE��n�=���=!p�;(��Zd�=�'�=�Y���X�r����/>�<�iD:��R=ֹ%�,���{�͇ἇ7<I*��o�<
%=\+�zݓ�E����>�<rK�<OԔ�]�= =bt�O9{�"nl=Հ�=�`�	��=u0�=(	��CpN=m3.��ua��Gﻐ����x���U:չ�<�>�~>	��ޞ�=� /=j���򥏽���<i9�@���A'�<H��=,w���
���ֽk%�=�h�<�����z�+�D���5��a4=u6>蜊�(W�=%��=�A�=�$3=�n�ڼ0=����)"�:o���̼��<��e��_�=�%<K�->�!>�Y���<�/�=�<t=�=Q1W��͐=_{�<KS�n
��Z�=�u��R3���ϱ<����y�|=�:l�ߪ��{�=Oĵ�����I=��z��(>z����#>H=[��=>ǎ:��=�⼠�=��=ゼ�����<V��В�<8��=/ީ���=�����=��=6<>\_=b%�;E
B��Ql=�J�=a}S<�ET�G��5|<����A�;�|�=;��<����ԩ	=p�н;�3>;:�=�޽��>�<3��=��t���%�����6�ܡ����ƽ2�S���u��AN�k�׼9������=䐻�
d�wK<�����=H7;�[Y=���=�"��Qȼ=���3�G�[=Arڽ {�<��c:��<�M�=b���>�=`TV��3=�G=W�G=S=���s7�=�J���0�;�W5;�~輧v�����;3�`�=v'�=
U�<h��;~���.p2���P<*��[!�;c��,�Q�����z=����;�F=�Z =��g={tԽg�S�{/r�����<=$8>���c�=˄��kg�=;����͠��w2���n=Չ�=~��yL�=�d��u�̽��@�%=/�=]��	�
>���������+�bi>=S_�1�&�:t�76�<�X��Ľ!�6a�V��<�˼�"�=���=�2�=p��=�2�G
)= �=sw=�[='�<tj�{���e�=�0�<�,X����{�3��=Uت�\�ý��=��7��^�=�S����Ӑ�<m�c�Ct#���6=����0B<#F<ž��5f���1�Ҽ�v6;�ㅻ�����yܽ���Xؼ'���d�=A�c=x�K]�p�k=zc���s$=��<�r��@�F=�Q��F�=X�<�`=��织�-<Ri�:V����=��=�U��9�ν�y���tz�=l���g���8��ҀA���U��<��f=��f<t>�=��1<�Ip�x�c=d�I<����`=*4�=��>�>½|�佾��
�����f<��1���=� �����=Sj�=e	>�H=E8�<�>'</>�������;/-}��ݨ=:_=��=r��="m0>Li*���8߽�8����=�;߼�=��*$>��q��s�r�5>����>���=�(t=\�j�͕��(s`�����q=I�`<����u�=C��=X>�R'�c׽�E�=�M�m-/=[N�=/�2��A�=1��;��<�����,\=]|�ڎ@�:������I!����=[�M����<����n���V�ǽ�ۖ=��d�#��<b�9�x��=u�<�7�=Ͻ���%�=X�K=���=[cr=eHq�����u��=.�`���<�*���Z�;-���B=���=vz�=	�Z=sB�=���'^�w{���˽����;���=��N<���1c���>�;��d���c(���N����
<�`��N���|�L�o�۫i<#�=`$9=��J=9=����T�$a��b��<'ǒ=Q�Z�Oﴼ�L�=t����U�=�y�<����Ĕ���#��I�<�=��=XU�ps>�B����=�s>�;4>2��|s�ԃ	=?n��dֽ��O<[�=��8/�"+�������xv=ʦ=� ����c=�=��<�w~=�����
�=��=I0==�e�+<߫��O�=q���νw��<*_�=���=����p=:ӗ�Ҙ��n��=���;J]=;1�&���1ӽ�=�s�<fO-���f��=� �Vs�;í�� �=l}���%=��
����=a.#=�E��9#=^H<�x̼��ҽ菞��,=%�=Ƙ����z; Kƻ�:�<g�����x�Ů�=�w:���<�1�<���<bn�=�U�=į9��>��=����1
s<�0=(<}��=�c�=V7>3'��z�9=�}�H(<("�\!��!�<�D"�A�>�|2=��>��=��>eĆ�zݻ=!"�=Ȱy=I�;;-�=�G�����E3��gǽ���:�����_�<}m׽�=(���>��<�x��'��B�=J��=+�=�C�=
⤼�^��[��"�G=�H�=}�=;���W��<��5=G�>1὿���c�ѽ��>�=����0O�<�K�<�c=�7�=��
����=�|�<�%t�_&=�w����EN�^J>x�j<���0���`x>f�4��T�ͅ�Ֆ��%m=��w=�y�-Se�POB:�b�޵�<ᑟ=/`�v+O�U�d����;ѳr�8F�=U�=�mQ��U<�?��t=7N���{����=;�<��ܽ6>u|�a�l�X&V<!l�<� �:�O=�1����(V���� >�%�=�^Z<�+= =���=�>�d*����<$.�<\�ּ��B���P>m�&��=�9�=�RD="Ŀ�
��=�Ȣ���9�[:�tq�3s��O�=u��=�>�$�2L�:��t��D�� v=�2=M,ػ� ���z�=��=�6����=Ñ�ߨ�z�����=�p2=�.�n�ٽ��=ϕ��r�k�Z?�;���u7�=�a���W�=f�9=�eV��B����=f�<���R���0���=�O�'��*�ʽ�Z�=����ҽW'�:��^=��=�`�L�����X=K�ؼ�q �d� ��;���c=�A�St�J��KI���C=�c�.j�=�Q&=e�>��Ƚl[ݼ�>�=b'�<�=��<����\�m��⼋ս���m<e�=&R��A��<f-1=2)�=���=������R �=��<=,��#L=�\���e��!�L���7(W�ö�<]�=����<ȂI<��=� ��>;��6��$�<5g����=�2��x��;:T�z=	Z��(>ZZ��+��=�h<v�Ƽ����඼��9=�ͼ8xk���	>���K����)���5�;����O����=}Ų��o�<���=�K�;ih��6ӛ��Y(��7�=t<=ŏ= �=�� =ʷ��t�d=a$ݽyx���G�=�"�=��>�b�	�>zs׽ x=g&�<@��=�C�=���=x"��Hn=X0�����<w$�;��$��.�~{ �̉�I+�=����ߎ6=�y��n�l��E�<��L=4�ڽC���C�J�[��/>�5�p�9њ=�mo<dK<�_ɼ�4��L6�,,<��	��|�<$I��EER�HJ����=e�R���/�'�ʽ�iH=ѡ��M��=��<U�;v�I���*=�Ձ��s�����ʩ<���<*����Ht�6��=w�v:=���x�'=F:�=� �߀:=��m<���=*��=V53>��T�"gj���= ��hb4>4�<�Q�<M�<>�ڽ@�0����<�3��uk>u[O��Ϥ=;d��6=5y��.�ȼ#R>�yl;��=E�=����:�<��=*(�<F�'<<]�<����>+�ݽ�{�=�-=���=�=��>p��=�ހ<�#���㽶�W�=�=�m����]=��d<��=i�n��At���-<z�ؼ�E<ۏ���3����:V~G<;����1�����<KxD�+tF�LqD=mƽ��[�(; �	�}�ֽ�a�=�5��B��6��=c�̽�,�KX��W&�=|F�<�
�Ll�<h� >�s�=$:���o߽�a�<�ܽ�1\=	v޽(���ʿ;���=H;����_=�E�=D<�=�~����=��׽���=�~��Q1>���V�<?h��-p	�A�N�F�!�f��=��~=�4{��. >2,/=�B	<X=!M����m����=�V*>��=G�*<nL>y�L;Ӳ��ߟ~;p!<7K���˞=9������W=�z�<K���ѕ�<�����R6=gPB�A�ܼ��Ľ��Ǽ9�/�-d뽢�^=�5=�Jy9�����1�]�<�%��U:��)>���<��~�O���>�2,����= ��;��;W�D��+ɼ�L<eפ�Ǖ=H���N�����f�����=�%*�`��=@�V�j��=)�u���Dͽ7����j���u�;�=]�ͼٜ��%T>=�쩼���>m|�;s¼�Qj=�����<x���ּզ��R^�MC	;�B�=R].�?̼��S�2�<�`=��}�`2�bί��ȶ����<�W�����=���<��=���=�>}=�-�;����/��=�})=��	>�]�|'�=�=��ؽ�*�<XÔ<o��=Z7��y�<<�V��cٻL��=�y<��=u���-�4=W�c=n�<=@�^=��*�Z
���ݽ���=�`�=�Z�;,e5<΀Ž�7�����;��>�$=c.滼�{=��=�`��s��<[߆�Ea��{��l�=e�=�w#>{��=�>l�>%2���"<�G==9�
=���=F~��--:��K��&ʽ�6��Q:>��E��!�;�/����<8���t4*=��м�Q=6]���t����<|���_;�=j��=�%��������/(�=;�g��r�=�o=t�=u5
����<lw�<a���q��3�
>Ε�<�=��S�=�����;2;����+>�[I�<.�=��d=gy =��<Æ=n����>M�=f��;AG�=����ʼ!�=� ��%=�'=Ѕ���ʰ�D߽����`I<���=t�=�م�0S�<�-½�^f�����L�0�v=%<��I~=�йtK���X)=� �=jE�;Ɏ׽��>�`�=	k��5>��<�s���$�<�C����;�u½�5�={�ν[Yw�sQ�=݆��! >�9�@�=��1��䧼bh� ������=�&>��)=𪎽���݆H�^r����=x8�=,c�;��=�A(��f�=�P��=I���=�W=��/�{��=BuW�6�w<��=�a��l�<� �:t]���T���|�=����5Z<=��>����Խ���Ϝ<nl��������UU���a���=�Z�=������=�*���=��i�Q/������C?<R�L<�(�fC�=8O=�����1>��=�K=�b=��7=��W� >.2=p#�b��=Q����۽Ƹ�;��=�V'��İ�1�t�;NK=c?ܼv�`=G2�<�L��p��%N�Y�:��ç�F�+�}�����<�<��L�޼�8e�x��=@)<>�M<�,'>c�*=x�����)=2�
>'������~ h�`��=<�)=ֈ���d<�g)=��=���*� �"��=M�E�6�=l>2;���=���=*�"��f�����<��"=���%�[�=�`�_�'��=u� �WU5;?©<6E�=����;=氱=��<j*�<*f��dhٺ��t=)�9=��ҽ��ݼ��&	���j��47�w��=�߽��e�(������F� b��P�<�c�=��d=�G���~�$ �<f�=��ƽe�2��<G=s�޼oK>��!<�5����<��=�9�<ė$>��=���l,���ѽ�f��,D�&���$���,h:j]�=;4=�,>%�Z� pl��4���:�=�P1>��C<S��=oMC>��G=b�=	t���.�<H,�=����<>U�D���� �<����2.V�AO =t����<0��JU���^=�З=,�g=��=*�}=�*>ԍ&<g�ǽۄ޽�<��>d�������	��y|=�9��JY��̬�� F�=�� >���tX�����<@>*��=��=Y|���=,	˼��V=�@��a��<P�=$��=x�=ch�<��n�bĻ��v=�+�=#��=�9��eƼD�������"���=��==��<��<���;��ż�����H�Z��=;�y=#Z$��q[�2�J����<��`���ҽ�.�="L�=u���푼&�>�x����=&��+>��=*K>�)����*R�=c�/<b��#Z��� =�L�<�"�n�<�0= 	�=�6��Zo=�{����ݽpy���r�=����լ=<dUi��@=�nh��N���ڽ�\�=����P��\��EC���S=m�f��xL=���=1�y���ֽ�r=BL=��ֽ�6?�J�=u.>	�*>S@=�=�^�wB����m=��<������� K��{�t<J��=�Tz�Ԛ��~J� (ռl瑽�Hk=�
(�Dm=�%�<Av�<A�b�>`t6��e˺=8ƽ<�S<��4��|�U�>|B)�a�2>�o���f��n�>&��=,%����ý�q�=Bf�^'O����=��X�8=�E>�>3P;v��=�r+=��<Y�{��қ=�7=���=��B;���;r����-=��}�<I`��j�`=�Eh=:$<��=/>�z9�=��E��/�P��PB�=�� >��<�=�v�����=�>��T"�=�k)>�J����e#=��=�M<>�=�3=�۽L��;�{��E9�D�=d��=�3�I���[�=|�=�M��ǆ=m�x�p�;�.>��=3��;����g,��m�<'%彬0Ѽ��>���=t遽��=�Z=XU��x�=�O��V˽=<%=wA<=��)����t���,��� ��]y������̚�|������E���:V��膽;�=��g=��=��<	eͽ�[�:C��/^��&����=c�½(��=�JǼ�)��l켶�����x���<�f�=9I7�	~���!v�� �=H�ƽ�a>���=�ߒ��/=� ��҄=s��=	�ֽ�����i�=t�뻔΃<�W����=�갽�=¢�=4�=��2= ��5���W{�m�ս}-�
%C��v =G	y���k�FF1=Թ�NU�<"��<�޼�����`��ΰ<�=K0�=�W�8�1��>h=d{̽�~���wO=$Î��@�<q�x;�>��΁&=�C�����{ۼ���=ʒ���<=/��;/�<��<Ș[��r=Ҟ�<���S��<�6�;@�%���ڽ �<B�k���;#³=ۍ�<��;=���,aݽy�=P�J=�L߽?]L�&����@V��׈=]/��f�=�� <5�~D=�(�<r�<j�>vN�=S��=���=�2�=�=�,D�@�`��ѵ=WT�+ti=�d_<���=N��< �_=������r�{��=��x=��U=�׼l��;��ݻ
�����,��cQ=��z���v��v<<�m�=�kĽ>7mn=f�<�p�=�N��t�4b�=�p�<���p�3��q̼�5���z=�|_=�h
�>���y�=o&5�0=������M��$�����c³��\<>��=)*�=FЅ�v-�<�.�=���=�c�=��=�Vy�L'�<w���cF��iֽ��g���B�Dw�=����S��G2�O����ؼ$e�]�2=�5�:�}�k��:+�w<�9����)��&�=���n�=�?<m�轨�.�{$ӽ�$>��=K>��ͅ=��q=��Z=Ս�<`��<���=��'=�0<�@��#��R�<>Zz���>���) >o^=&��X>�0˽h'�=�`=-&|=O��=���=G.=A�V�ŇJ=�Ȥ��ū<���=��K�OHY�kxC=$?=6��eD>�s�=cQ��a6�H�� vƼ��*�s;e>=qΞ=���<�/=�$���=�V�<t���4;S2�=4��==^8�7��'�=N�x�'�=��C�>��¨�<$98=Y�=4��=���<�4�<r<���s�=�k=��!�L�N��=�`��n՟=�.:��ب�e��=`pý�0J="�ϼ���jp��'����@����S�>�o���>)��=݄��nhý���4hy���z�W=���Ț<�)�=
l3�B2�=*	��Ǽ2�����H=h�˼�x<=#=��߼qA�AU
��۽?rZ=�0�0�=��=-��n���R��$���V��=F7=�'R���>��=��G<�y\=�i�=�U�<9�D<�CP;3�k�񬋽��;;��=�?�<5B��s��=_a\����<DL�<����/��ڭ<=���;$x�<F&�=*�����R=�˫=Yu*��I6>��=J�B<��ȼ�1P�S�=��="�b=�/���
��9UG=6�=�J��[���X4�x8�1����Ӯ=����h
&>K��<(J�=J��<T���35Y=_ݗ��8�:�cn�t�)��r>�)q=�d^<1a�z���PT_=��z��L=��Vӽaz�=g��=>�|=��¼d��=_ ݻ�@}<�ے�����3 �<C��=��\<�o�=1��=<;@=� F<��<;���ʠ�=��Z<�>�/�<�ߣ�NI���J�<��n=T�üJ�x���k<c�<��^��-��?+:�O����=>�5> �J<Қ�<� ><���=��=grs={��Ɨ�BᎽm�=���I�K��8�����=���=I�?<��R�3�u�|�=�LU��<Z��=Oކ��T�=6#�<�M���>�
V�|
��M�:��\<-×�*F<=�~�t=��>���;�'>�	�=8<y���k���Ժri%�녜�EKM=�D=} X=������<�`��&�:>����?��;@�W;�L>�!���*c=����<�<��;��;PR���B�x�Y;K}�r����ˊ��ﹼ�7�=��1=R��=q�F=��'>��<���<ߌ=
Xg<*m�=��������<0c��_��=��==��h��=�=pM����¶ >xy��+sC�	�������N+���7����< ZE=�dV���<N1>v,���Ѵ�
ԣ<�@�=*Fi�q��潒it=�t=�7�<�p@=Vap��vP=�$d�%��;w	��+Q�=�qI�-��=��=�C�=��=�� �|��=C�;1�=�3l=�����	~<o��=��n=��Y�܂>�5=�|�:μH �=S�=Z>�� ���<B�r=h=tw�=?�<���=[+S�ݎ���y������)�<�X�=h��=������<'��<���=��=����?�=I�=J f;y�<��;�+���It��N���S7>���]n۽o^����<�)=%�=zĳ<B]�=b9�y������Ij=���na���y�)��=��A���l��R��6�����[8o=�Y�=��Ž��=Z�>b����+�<�گ=��	��Ľ6�<�^�~�G=~R=��������=�7t=9bŽ�:�w�$<�w��W"����|L�r��������>�
=���=�&�AJ*=[V=n�T){�y�� =���e="�u���E=�$���?N�@��ζ�=�㩽�#�p
�0����;<�ZW�vy��"Sͼ|F��uʼW����7#:�0.=-����\@��<��<�ý��|=o� �U��󮽦K0=�M��s=���h\4<��/=����/���
�=%�=�e�ӛ��Z�	��.��좽���<ART=n�V��z�=��{�y/�<�&��-��<����H�7<���<��d�?�;.ͺc��Z�l�q�S=�I���[���_���4�w=�M���=ef�;��>�˒<�(�@&d<�ͽ=��=�E����=�����Z�=B
�� �^=Y�3�f0�=Q��=A�a=�Y>i�7;`�%<����	Ἧ�x<aH���<JNI=^�Z��<�E�<��F�ս3�}�.��� =98L�D��{���>����7����=�
<�Uƽ�9߽%я���+=��v=�Z=t��=�S�_#>���=3���6��<|n�=g���[<n*Ƚ��v�t᷽�Q�=��=��=(A��~���G	��8ּ�R=��̽�H�;�E-�0�~�==9t�=�*�=��	=��=\&�< �z=@-�;���7�*=u��: y<��==s1����=	�`=�����<�=-���O�"=$�=�q��=0��<�\��w��м�"�=��=�����h&<ϣ���=�=my������+�=h�>te��e,�=��=�G'<a}\=d�= 	>�~�����<� �ک�=^���3�A=#=���;g>�|�<􂮽=~}=7$+��#�<�۽'�b=4\üks��6
0�o��=`�>�>�=,�/:R��<������=\׳=��S����>h��f�6=���߿�=�Q��nٽqdC=��=���;=E���I���K.�c+>��=m:�Y���i�|@���{g�=��Z��a4�����`�鼛-�=�м�n��	}ļ�<�=q�B=�AM��a(��-t=���=��>;b�f;����Mk=99?����=��;Oy��4��z�j:V�5<���uZ,��>�=�e�9;3-<M�a=F�I����=�E
����<���T���-�=�䈻-o]=I���=�Kd�����Q�P�=�M���d=�?�=�8����u>���� ��>�>���;����}�<�� =�=�M�=ص��(|��|]�;=z�=,�������x罞4��+�=��ͽv��0=�;F�>?ԙ���*=x�����=��>I�=��j=a.n���	����;<�G���=��ν{m2<�#�<���ꍹe�A�4t:>C�=��V=SlK<���<����Y�9��8�=�v �}L#��r�;��W��m&=�;1=:�<�9>e̽��=�)�[=�����_�����?录���>T��{Y�?i��G�=��=�E�=1>�"�;#!=��b<�r=�7<-�����<�t޼!�����;�dý���=u�=��'�u<8<�5<����Q=*�=/n>�=I�<�=�]+�Ù�=þ�����ܽ�N�l�۶l=�Q�=��%����=$W��4��<�� �r%��ߺ!K^�y����<��!<�	�;�[R����<f�=45���e�<թ����<��ݽ6�=�؋��O=�����V�=3��=��7>��)�N�V�bB�@��;���=��<���R����Y<��=�_+���A�����,*���/��;1+�0莽:��<@;e=uUC�.�>5�ٽ
G�=��h=�1ݼ^��=pؽU�+����<^�=�ʢ���S>��<<[\�ڔ�����,=�1��6j�q�����X�6P ��Y��s<*(�=Ír<M��*�;Ͻ<����\W�="�={������R>����V><R¼m/9�`��ٞ={�<��Խ��g��#;�=�3Ƽd����>t�>�<����Z=<�?�=se��\(/��g\<�`=OEp=�K����､ϒ���=����-�`�O�����	�>���A��=�ʲ�s���>y�<�}�S�l��E= i=K��$��<5?��x����l�=�V�; �=v6ٽD��=�i��#<�/*��W�<��=x!=�>cbļ��'�
伶ky=l�6�%�<&K�=�uؼr:��u�8;�\B��v轏��<���CH�i���ƭ�Ε�=�����<ߧ >|��mz='E!�����2Լ̾�;�;�=�ؽ^��=&��.	|=�@����=�rm��]�<���<����nJ<��#Q���<۹=&�=�}ܽ�М<�'<QW�<��[�#�<�˼W$��T<a"�=��ýN,4�ԕɽ�$�=?c���;���9s埼�6O<��s�j==�B���ę�6R�����>����o=s	��g��Gc>�Bq=�,t=�>����<7��=���=����*�������o=I��="�]:\��;�r���r��x���l�Ƽ��=C	>cݿ<���=���ɿ��z��:�����ڭ��﫽�����2�;���=�<�ai���E�ʵ5����=N��.NH==�!�*�L=���L���֜G<��齣��<������=4��<��>�H�={}��q���!��_��<_i��.�>!5ݽ*vX=[C!>d�B��P��F��=�_�:t1�=��ӽ�?�<�/��r�=b��{+�[v���ɼ�PQ�X�>� >�+=���𽻭���)�������H�=l*>]b=j̡����P)=�.{��ኽ�,M���=�	��+���p
���ɽܟ;D=�OE�s]z=Bqb��
����� +�<,L">�爽O��39����<�$˼pm@�J
<Q쯽)Y�����G�<��(=���[n�;�4���d�>r�[=��Z�9[�_�����5�ͽ�Kk����=��ɽ�q=����!\�jM�;�f���j�D�T�ơ:����<����*\D�H�L=�uɽ�=m�=y�z�������Y��nQ��6)� ���;
2�=�1�B�=��=^�=I_�cŉ��z=&���-��<�=����X{:� ���K=�ύ����=���<��=x�1>���[�=�h�=d�>��a�}26<x���AK��Z�s�=�f �7Z��z$=}�1���=��Ѽ�����v=H �Q	��$���~�Y(�=\ ��ӕ�>��<��_��-��N�=���<�m��_�<(�=ͅڽO
s<�CǺT���)!�=�W=��c<��>��I۽k�ܽq�ɼ��9�eR��=>(�=���СS��R;a�U�G}=���=�#=��/>��)�؛l�`k���>���y=�ђ=�����］��=��=���4�k���=d;B<�������s�h��;8-�F��<�3�G�<-���� ���d����=��=ҿ=�Vz�=K�w=��>����[ټX��vח��ս���t��:�=p]�����v��Ո=�P���=�k�<��>�Y=$z�=7p��$�;<Կ~��'P<��l�
A=�d>������< ��=�n�:m+�;���t��<[�:) �;IA��-{=0��;�DX;QS����Խ��4B��"�;������<K]>��=�=�=��p=Իٻ�����<�z��S6���e�=��;���aԉ�� �T�:�u���j >���M��=���;� >���`���㹽�g��<ҝ���<F-��Ǚ�>d���>"+�=B�!���G= |�=��=�k�<�&>V�t<|���C);�*�(�Ԟ<�b$>�kZ=���v>��sR����<�w���G<��5>+<�OD����=f�C;��������<zl>�ˡ���=N��<|�E:Z\��pu�;cv�<$�=��7�z�A�=�i��yw�=��=O�=����T����������0��.��;K��;���oQ�<�K=o�	�ؔ7<ҝ����W<�c������-�۽yǽ���=��&=zE�Z�Q=/��`c=S����掽kR��콨_�4��J$�Wuؽ��T<U�A��� �GN�a7Q=7�<�D�;����D����<]�=ұ=��ӽ﹫���ӻ}��=� ���=^I>��<�J*=C��="��<V�����yS=)m>�P<-)ؽ�;�;�;�a������,yf<[�E=aA<��S=���=�O�=�<��~�l~����=i.:�g=�,)��p>"&�<?x�<�C���0���E�=��z=�)��,1@�Э�=�i���R[<�G�:ʏ9<�R����+<>d�'�t+�<)��Ʃ�;iE�==$�<���}������=L�=c��$H=��N=]z6=�Z0=���:x�x�O���~=A��=��ͽ�9�=m\��C<w�>�R�;�L�='����Y�=r\=�d�<A_K=l��=5s�=���=�t��au=��)>��=�,���׽H<���+<��;q��=��=��ټl�ؼ�3ὐ�s�f��=�mu����=���d�#=��ཡٚ�N��a�J<)⼶z*=8N�j�L�e�>�ꅽ;��\ֽ2��=��=�4���t��񼴽��߬=Xf�=�l��3O<���i�&�c�J��"f�=�׽�7w�=�����%�"�xb�����/v�=i�`=ϭ��qD=������'=��= �M=󃝽�w<i��IP:���<�)���=
�{�N��H��$<ü<�~=\���Ƴl=o�{<��=@G=�ki����ZQ\<W	�[��C��S#�D󽫵�<�z;����=+�>'=�q����	��m#��X�2zx=T��=0���XF<��>\<�9<�����nɚ��>��=�E�=.3�;c��<�����F=��:�m<�)�:�2���-�|�	�����EcҼ��K<	�>kM>N�:'w�hi��uP�=�+�=�>2�ʽ��?��I�����=1�=g\�=�Kb=��=���%z)=+ǖ���=;ym�)W	>����s���,�����s��nAo�	0<��1;�3�72;.�<�x����=:=�K�=���=��<��(�Ea׽���L��;��=9c����T��V�c�����N��B����,=Sð�W��<ch�3�6���{�V�S=�'&���=��h=��y<��J��"�;x����5>������:᨞<��r��A��Ȓ=��<����`l�=G��<q	=��?��kc�������[�]����8D=]$=�V��{�=Q2�;�ݍ=�=�����9&�=�>o��K�<O����N=��&>��½��=�<x��=�1�=�B�<�`�=�\���o��T#=�5W={�Լ���*bѼ:"�����=�� >��=�L�<h:�=�Y9�a�<�f�m����.>��҃�����;�=���=�^G=���<������C�=�&����)=�v%�y��=�s�TE]< �=����y��;!���i/=��ʼ>�u;��U<�~�=�p���=#�<�!ϼ�.-��ȼޤ��� F�7�
>H���&#\=^Ѣ�c�_�K�0�.>g���h�k1��4���dK=��<m���;�= (e9���������<.锻?�-=m�<��@��u�<g��9�=� �Yi*�'?ڽ8�:��!�=�]=������=�`=/s�=4�=e��=0���
����B>2�G�g�:��1�Z�&>tL<�= =Dm����U=�(=��=��=�ݯ�[�-=.ț������D=̚�+ݽ�$�=���	�����#=���=P����Y=3惽G��TB����K���S��K�=�Ĥ=P��=�8��*�8<\=���=j-ܽ窙���<�4��q�<���<��>1�v�����f<a��=���=B�4=}&�~���bE��kY�c����.?=��Ὅ�f���; ��#��M\=@M�����=�=m;Ѽ��Q���>�%�ӊr=�F�𣏕�S��=ϔ<���;2����=IK?�m*=��>�)=ĩ�=� �m,L;�	����B.,���ʽ_|�=��=� ��<�B=�餽�x�=g8�=g!�����������=���<����G~�����Xt��P7�c�=V�d������=N� >��۽�U�<r��
�]���=]_�"���Z���{P�;�穽KiK<�T&>(u���0^<���=��g�`�"�{��=�r���m�;�ԑ�9>p��p���i=��=d��<��=�H����=��ὸ��=,��<Z>������~�<�8v=�a����u��=�:D�t�=ڒ�^�=S���u���vW<��;��v=�*v<��y�Z��&n�= ,���^�=�l��3�[���!=B�;�I����Nl<�#�$�=A��=E�=�-;���<�?���=���=^��=v�7��n���A8����Z�<5�l�K�O���=sו=��:<Ɇ�<P=��=0�K=�G�<�l�=j4=��;���1�z��Z<��W<���N����=�W�<e�,�[k�]?s=���[��N��,=Ͻq�=q�Y��#��z��<W�;d�����=�=������,;L
�<6S�=CI��I�콆ұ�μ��=��
���6k<�2q�|�H=d��<�>T]<P&6=t��=������;���<M��$��=~��=��=q��=,�=���<�=���>v�<io��	� =�T�=�� ��#߽\%"�ī���=���=36�<8�üj�F���x�`*�=[#��Ld����%<T�AN����B�D�	�S��=���4h½�g�0ξ=�}�=oG;;r>L��=��\�H�L����e�=�����o�����<��0�E8����=u�޽�"/�2z�<A=쟱=V��>?eD=]�<�EF�z-���a�h�&=�ͺ=�s�����<}����с�D����:	t>zIN<���� �=cy����hq�N� �(⼻�k�3i��6�;~�@�;��<�=ক=ԛ>.c�a,��JӜ<����߇����>=��V=� y=;J>�l�;i����9<���m����=Z�M��hh=g��=3VD=��Y=�Z=!Wu�:���zF��e���E���E�����=�H�<���=Je<�i�=�#��*�=��߻
yt��󱽵���q��Pb<�j�l�'���o�Jk���:�9&>���C���8n��9��Æ�<s$m<OeżA��� �ܽ`Y>���=AR
�W;�=�bd<���=aP��L�8m㺽B�=G.��H�=��>n�P�`��=����SV��� >S�*��Nm�@�=Z4���k��� ;��ƽ�Z����=T�q��b�=\�Q<��=s��G��=D>+��=�2
�o\�=�+�=ԙ�<s�!=�N��,��ќ=�����)����rZ�r�:�]�;ʴ�=#�_=�춽:뽑�,=ӣ���\g�q��=���?�<p>���=Y��=�7> �Ľ~aͼ��;d���E���A >�ֳ;$>���<YѼ�޺=$ >�^6<(�;�7�=�w,=��= x��Þ<��I=/*,�,�=e��=�k�<.J{�\μ��~�<���� �=��=�V]��+乭 4��e��ž�:f�>H|�����<�<��=����{<�=6��<��Ȼ���=5�g�ķ��P"۽@�����_=g�S�x{�=�b���b�<�b�=
�M����0䑽F3�����y�]��YV��Q�=l��=R�W=�5<i�����>�e�;�:`=-�>��=&�p=p�Z�W��=���=�8L=�1�=���=b�@��y�����<�?R=�n��>��>�W���g��є�<]��V4�=��=joS=�8:g3>�>s_�;P2�(�Q�bƷ=��E�X1=�ψ��δ�99�:��:�쭿�����+D�p�Ǽ���<��"��X�d"���$�=-ٻ���M�����|u>����򉂽!�f=�>�<��;��=k��=��==&�=�I=����������\�Û�;xyQ��n<���<�a�<��"�y8=Bi=�:?���v�ȧ�<���������B�F=G�=���ݩ�����:\���λ�Žy�pH�<+��Z�f="�z=��=A�ݽD{:���ʳ��F󔺼q��]0��T=N�<^d��S�=��</���������!�^��q���-���n�=����(?�!G=k!"<�8 ���T<?L��訋=�r�!�$�Y^8���0��x��Qbv��$�=����>��ռ����J��n�<t�=H�J<T��;T�=�t�=�jr;ս�؟=ǽ�������= �f�Sw$=9�����k=9Gk����i��=`�޻$�=�c=׳�=�h<��(i=��<�_���]��r��K�ŽF���:��0�=p��;8�=PL�^=�ۤ�"��=�c����=n�"=�ʽw�ļ�5�������׺ހ�=nm�=������>�����m=�h��T�������B�=YϞ=nA =f৻fk����R=��缮s��W�=�Ts���S=F������=\g$�gS½ŸM=�^�����;lO��O#�=���0>��&���P��<�*�=���< ���o~���i�=�ا�
�O=B�=M��H�8�U�S�2!>���7���=������=\�ϼe��=�_=�F��3�����=KĲ<Z�{�Nv��T�6=U�~=K�={�q�����ϑ˽g�=m⌽�b��6I�����=hF�s& ���=�! =n�引�̻ë<�K�=ĺ�=��	�=φ��[ ü�.�<��>иս�q��w�=Nd4�v�<�	�=�I�<13�=��>����]U=V��:������X=ȗ=�l�=L���nՖ�8i:>�ڻ=�O���ɽ�rU�B�=�6�=;�������$ ���;� J�㆚=7��<u=Λ��7[<M��ۮ<j����<��7�n,�<ڮ �q>�<ӌ���ٍ=~���Ί>8��=Ϸ
����<:>H��T4;t	���ﻖy��~�澪;ٽ�)�}�{����=������bn��S����������f����-��=��d=��+�gG)�tӭ=Iμ �G<��>��<���_�޽��=�yF�e�Ľ��=2�=��>=�\d��^C<�����<;����L==��=����c�s<�>�=��<�ɏ=z�s�][�<�`�=;9��Z = ���U8�~~�*��:?�k=Ћ��֣=���1#=ï=����u�=@�=�&�<k+���g
<�3��V�3�k�{��h��	>3�>�$��<�_�=u�=5�=���=P�=P>'@1=^��=b��;��!=a�>�;�=���<����h=�A�=�kd�����{�����g=����$򓽶�3���>���*�W顽�?鼷�i<d=a<nK<�,�(���4ݢ����S��<�O;^Qu�$�X���=w�ѽ̓f=���o ��F�1=5���ur�=���(��k��;t=_���L=o4�=6'��5����=im���s�"q"���Iʽp�M�<��=FMϼR�s<�r]=q�>�����D<=ѽ���ȋ�!�Խ
�"�ҞȽ���=�:�;<�<�~���Ƚ�8�=4�G='#��E^=ھ�������˽�q�!J~=�Y���i=g)��4��g�<���
�>3�<x��<��ռ^����;�]��a,2<(�>T�
=��8=7;޽��?>���P�G�>4���n㼕��#?�}�8�w���ty�F�G�=F�=K��� Y��s4T<z����N�=���+M��Vu�(j=�3O��5�<�H�=��<q��X�<��
�0<�Z"�_C��{p� ����R��U����<ԟJ�����<�M=��,���>=)����w���>�����%�=����9��<v����ί��݌<�����=��>�XK=��<���=���ĵ�����
!���B;�vĻ�a��B=>��=<��<ĲŽ0Q	>z?�<� �%׽(�"=Kn޼5�y�I�B�4i���/��w��l==Z>���=�w�=Hޒ=���=EG�<��!��<������<=���=���<4]=�$�W�g=�#�=r*���<���u^��>�<���=bL=�ျ}'4�x=�J0�ʲ ��%>z�P����-TY���(=>�>G=�R>t�G=�c���=�?���+=z�y�k��=��ɻj&i;
�=�1��q:��o��O���:��Չ�<*�\=�:�=/�T�=k�=��=�E��\5(;��˽N&���	�@U�=c�=o]�i�=������#=m���+ݼ_�>qs.�&�W��!�8��=|>��Cdt=M܎��j-��=�h5=�D=�.=<�L=�^⼦>P�3�򻨽#����]=dǙ���;<�v*=W%�<!�U=���<Gb�=sMȽ?���(�t�ͼO�h=a��� �-=��<)qw��V�@J��B=���=����^N=�W �w��A������s�=��y�G�Cr����Խ��9=�̡=^Ì=4�M=x��=r�Q��üD'������S��8u�蘺�+�N=>��<v�ϼ�bս�� �ҏj=��ԽpL>�m�=�b.;h��=hM �̼ͻ;�=P��=}T=�@�=��̽�廅���InI���%=T�Ź
=F�����@=)֓��X޼-	�������|���4> �$>���X	�1��=���w�;��+�U��<�l�=�sj=���=� ��=7?'<����_4�Ln�;�H��y==�r��S걼���=�����>��}�*H�@+=m��=k豼�fq=p�{<��_=S>M��$W����<Ho�<�o�<��>�E`<�^�=��=���=l�<���E����4='�+=����Q�L��Rh��,�=d�=�ς=E*��
>�>�?=�g>e�c=%-��q4=t��;b���D�=�� :$n<Nɕ��(5��Pv=	u�=_ڈ�@lǽo����J�*��=��=؞C�m�u=�q�[²�,�
�3�=�t�=�->|.>L:�����?c���,�<�F>G9a�N:�Hm�����=3�y=I�=��� �L��{]�WY�<*<7����T<O= v�<꽜4��^��<�w\=��e��?}��X�;A�ս�}��D�>8�=�PZ����=��=_!=A�V=�2�=P�̼���=|��<P1�<��=�Eڽ����u�B�U[�<��D=3w�<������ǽ��T=�v��W#�4���G��<OW�<ӑ==� �H6�=��=��ּco��0y=s�;���=��r�׻h����%	>v>xJ�<A O;%��=��
;֌�TI�=�؃�A��=�ļG�>�צ=](>G����I�=���;��b=ƴ_���R��nܼ��I<�e�="��Q?��fm����=LJa<l�p=��׼���=챨=^w =T�== ��=Y>x����*�=��^��Y.=?s=��<�=�t+=�;�����2{�)��;����^+�IO���;>>�=�°=�1�;�W=�N>=[�<�2��=(������8=5��=�׼�Y#<�ߪ�}ef=Qv�=ŞH�(��=�$@<�P >y >�K0<X4�=���!�=#ڻsv=��6yռ�}B�IB< �>>��9�l4��1Æ<ie��Ĺ����a`z����TL�=@/�;V���l���4`�.�!<�">t�=��;ޖ>�ok���C=�J�<k���*��=m^�=p+�=�`���t���	=����gu=�%�F�/>�U�=�[V=���=���<u���n�m&��l=@:�
��=&�=2�˽z�6<e�'��2��z�"������=ϵ�=��=(�Ѽ���=x�^�=xD;�K=X6�=��?�4�=)U=Qr�=�=h�!��I<��_f������Dڽ��h=�=�h��	�(>�ܼ�h�=8yQ=r~�<]�=�W@=�u'>�1>�� �ʮ�+*���2�=?^�=��2��@��w>B��j�/6�=��|��=j��;�/��L=ldH���>�2>��K<�=�,���i:]�=ü�􌽲0��XHҽ��:�hA�����=jg$����;���;�F�<�m��tr��t�+|�<j顽�><%�|=��0��|��$�:����R�S�9{��<ڼ���Љ-<zQ�= ����8�K� >�Ľ�H�=�fh:3�=�{�<�>@=>|�<&B��^�=�O�<Q�=L�1=��;:�@
=s�=��= M��MV�Fɼ�A=��B��]&����OB���j=#	>ğ���H=���2K>�b�:P��YH��>���<�t�<Rz��Ni޽�M"=�'�9��������+�n�>}�;�]�e8=I�ལU���ܽ��!>B������=�����=t'=� ����º�V��+�޼;��<ރN9A���q=+>����ǽ.4��ͺ��o,���<�/6<ݟ�=��<b�O;fu����_�<?+=��=*E=u��������=�d����<��8��*h��'"=V�>N��<Zw�=��>��=��=D��=؋����>�r;7Y?<M֋<�>�����k�&E�=nG8�;��bn�=�l��s�>I��K<�=�5V���9=zL��8M	<�X�=J��	�|��j��ǅ=�P�=gE^<7��<}惼R��<�a�=��d=Ur=��|��0@=��	���=ͪ��P�=��<��E�@�ü��P=�B�=��?����<��<�c�=x=)����C=bc��#���tP<-�C��$��j�;s�=��P�R��ǽK��<B<<CY�=>���>97��:��;�<�=圐=_Ʈ���x�`���BM>b��,�<�qn=���Pk=�CϽp��O�=V�=@=��N=���<��@��=�!>=�⭼.K~=!���{����>M���W��,��;T���*�`=�<(�V�=�k��+**<��s=�a�=@
�=�*�|nm<�T���=V%��q�n��;�F%%=�s!�$ԟ�e���:��~�=ز�=�=��
����J=�8V=��<�>�=��^�A����t`9���<*�׽
�=��N���伌)�=�ڻz�=h�R=�V�<]dP���~��#�=[����=K�`=���=�9.w���>	K���<:�=���=����
�u��xq=0�^=�.�=]��=iZ�N">���<S�����=t�t=������=k�i=֓Q����H<=$ӱ<X7>�Վ=B�=au�=t��=L(ƽ˦����@�f��<�=2=���ND��D��>�B�K��ڼ�b6� f=(�T;0��n�<
R�==���<E�.=�&L=s�޽t&>Q%>u�>DP�=�w!=c��<F�=� �=x	=��3=�K=�j=�q��9+�>Q	<��<�k�T����ک��yȽ��9=4�m�Ҹм���5�(����x�<t���e��=�c0=��=��I<��<��>|��=�5?�����p��r]�b踻?�v=`v�=2P�zwż��
�پ�-,����<�<�<���=����9�<+" >�h#��8=軝=�,�;L>��H�=����6S����y���(��ts�Ԕ���mh��7;�Fc=���<;��<U�ս���<߉�=��@=Ed8=pvH���b=Q>>���ߦ=�抽'��=q�ν(g�L2�<�����A�=���=5��^#�=.���V�"<��[ɼ=����H>�%���A�<�<�i�=�w%�&�>��<=��=u�[�d� �W�H��V�=rԒ<��>�"r���>[���m���x�޽rz��b���2=k~=u̼��>��=��=N��<�?!=[*�=;��=S�<g��=�w���O��E�=��,�����P;�q�=r��="2�������H��.=;���<x{4=�;�4�1�g���/�=��<�Y>�;м+a��z8�=)7����潂
�<�=�/�=�q,��/=�,�;�Q|���>�,�=3�x<ϰؽŀP�^�f=���=��a=T�g�W��,�<�f˺rB�<��"=�Q��u�8W.��l1=��C�&�q�����=��V�>�F=�/�<8߼j� =I��=��=W�=o�	=���=z�{=��r;D==j�R;@�y=�Rܼ�s�����<�a=�+�dIr��&�������"���o���<�>�/��1U�pc)=,��<��>,˔�M�������=`�l�%���vk=��<=��=$u��(�=Kpq�⚼��`���=�顼�=�:�<Ԫ�==���=6QO�/#�<�3!�����S;�q����R����r�</d#=���=ʬ�`�>j3�=:>�=�!���(?=�G�<a�=Oڼ0�<�ȹ<�~�;��8�)���=�?�Ĉý��#>	�<pʻ�DK&��*��6|�==�������=ُ˽I<e�G�,�2;[=B��=�^g��bü[�<M1��^Qƽyi�ـU=�q<8����=��=B��<:���=�q��T�<��M�B+_�}�|����=����cѤ;��E="S$�{�;��<1����=G>9�*>�c�= ��<a��bxd=��=�`�<��Q=�I;�����-�YY�:�=$3x;EM��<l@�XW�=Y��i�>��p=H]=�<
���[;�$�=�ͽ��>�i��C��=gcx;��=Q
�<��ȽJ��<'��<�!)>�Q����P<��h=�;<���=Ι+=<�V��49�ԏ<2c�����Mλ����J+ ��m�=��	=b��<��f=Nk	>G�/�j����<�����m̽�!�Щ�m�Լy@ʽ��<9Z�<y-�=�p>��=xx=V�乖}Q=���<p=6�6��["=zϽfr�=M@>Eؒ<�)<C��<��3=d��n�<�Ԙ=�����U)=�O2=!��[=(���=D\��%�=o���.=�S�;��(�cL�=A���`�E<z�̽a�v���<�;�����=�<�����ͩ<����}���5j�a���z�<%�>�F=�<��Rx�=�%���I\={Ľp��=��!=B��nN
;�ὑ=b=V1x<P�S;���FY%=���<�">��ֽ�s.>���=Ԟ3�X� =�^<=(Խ"yH�%'�=ғ�8��FT��B+�H=���@�k�j��g='�I=d�k�P�=xMU�ܼ>=��z�Gf(�Q��=��;>�h+=K��
� �;f��=�eR;�Hi�f���g��!{=�6�=�3�<F����K�=�p<���=,�=Ʈ��D��+'ǽy��<?�=6j�=@�<�駽��ջW�<De��3;T=1k	�Fڼ⣴</��b <x�<�r=C�$� �A�����<�u��f?�<pք<!N0>*e�3����[=�<�d�O���]�=�D
��f����ж����<�q�s >�Ƚ��=���d�Y��Y��8�����=��(=��v�.�=���=��=�uo=�N��=m=w�= P9V/0�0 ]��t�:��=2��=q*<>Ԋ޼��<BS;��,=i��=f���t�<�H�<�:��������<i�W�aF�Lp;졎=���]k<2�k=&_׼zL�I�7=��<���=rI>2�*=��=/���8t�cg�#^=���<�p=�E<:@!>��J�d�=�����<#|���x����^�<��<p��=��a=�<Ba#=}�;�3B���AϽ$��Q=�Z��~{�=��C���=���˚�	� >񑵼A��<^❽m[="N��S���q�<�D_<���=�F�=ۥ=X��=��>Z����=��>KP��E�<�1>W@o=^)
��&k=_ �����=�`����.�!U���� =V?�=9�����Y_>�N�<�<��h���<�s=�'ֽ3��<�2��V���V?�<ԿR=��&�0�Ž��&�늏��wY�~"��Q���օ=<�(�0�.��="�Լ9T>��;:�I��~ټ��:�P:b	<͐ɺ��t=Oh>����Yl=3<���>X�;}�q���нĽ�<U:�=Vg�4�0Z�f׊��ط=�F;�R!=���=�>���<����"��<{+�=�������.\�y|�=�1�<���=H��X��"WK=)��;���=��_<T�{�����A-<�&j����=�T���=(�ҽ��>��E
=�&��0r�=��=�M
<i�P����(��<�-M��=9됼aWh�d���y�=��߽��=�*<|@0<�!>���ӡ|�Hi�4�=IP�=ڊ�BP��5f��aP�=�)� �U<���+.����=wջ=�= k�=�7Z;�Ǆ=n��O�u<�?Y<c�<�t<�����/w��J�w�>����<H^�=5T>!=�'����=���5cν'�<x��R��P�=�]��>��=�&����NZ<tã=��D=��n<7]!>l��<N8�;b�V�	>qt�=�N�6y9>�%=<6]�_��;���J�<_���5�="V��5�n=M�-�E�����=�M��	���k���#�i���0�;�= #?�;���P���Լ/<�����<1�a�0t�=��l=���a�1=�@��Zi�����+#>L�'�0�>﬇:7�߽�H=C�><�g˽�&н�Z�<}��U/�<���!k=]
�0��:�=�;jу�=T~�� P=J\>H�=��������<�G	���9=h=9�i�`�z��bX=�v=�н���<�I��Vs���w=O����;Ӗ�=�j=[z�=b��<RqK�%�
�7�'��=��Q�ʎ=�y>�X=7�;䗜�}�=���E\�=t�<�䈽�}}������l=�_���T�;��a�~�v=�C���l�=�c��5k��b�=�e�<��,�Y��<�t=?�\<KO	�'��=g���=;'��4��SL��Yq*��w��ټ,h�<�>�;/� �(�Խ!|8�l��:σ�A��Nc<��꽝�=�+��-=O��
O="�=�y���}����H�=�:��>�=���<t����&�=�л�u��0�]�K�<��=��#���l�S�=7�"�L�=�
�;�3<�7=��p<�xM<d=~��=�	>h��	�u�Ƚ1?d<FmI<fj��lT=Ao3=�QI�k,�א��8+��Խ,��n�K������=T#�<E܍��ܜ�rV���ͣ=W��<�D���>�P����^���VŻn,���9�C1����;�J�<�Z��ϡ#�����1���1D�<V	�=~ꑽ�M���=0����=�����ӽ��=��|�N*=�yϽ��y=F��=�������n��<!�Q���#�<?�Y=�N =b5�j��Gө��$����i:�{�=���={T���5��ƍ���ҷ�R�N�R�[7����;������6�`$?��1��`���I9�P�b=\X�;�#���ͪ�~��=i>�T�=���=�I,=��O��<nR������>hMJ�[!L��p���=���$��<B�=c�ʽ�����=�L`<Vo"ֽM q��o>��:�[�=�4�="�
>��c�ҔͼB��<�p��'��=N2:<���ƈ��M3�[�=�ވ=�yd=��=(G��Ի��y�>�T9>�-.��4 =_�~�����x��<:߫��Z�d&j�H?�<
-;��ּ"Y����<�[�;��<c
�=�ۮ��ؗ;�i�=6d���+�<P=l���	%��~��rӽ�Ug=r�����<-@�=�=�;S0�� �<�c=��ɼ��=fق��6x=�Ӂ;�#�����p)/����;�%���C�����k��a䩼3ʔ� {=���u-�=�&9�������=��
=���=���=�ㅽMP\=��=�(��V.�PG)�Y��=���=�s-=Z���{�a�«�7�<`\���+=���=@!"�Ylt��F�<8�2;m�*<ճ�=Q놽7���u��;��
�b���<�g�=��/��96�'W=���<W�ͼ;�>����<�=t��;3Ad��S�=�s
=`������/��=������ѽn�=T�<i�<���􄙻���=؆=cz�=F]">0Q�=Sf��}=�ޫ��2�d�=�;f�c���h�=�.���뒼�$=I�^�Iu���b=C�
�����{;A��S�=
f�g�����<&�=������^=0;=`��p��;Q��=0Ȼ=t��=~w������ܘ=�/�=��7���=��>���T=��U��ҏ<<�=��x<��Ƽ�Q=J�Y�ۉ=��M��d����<�c�<�(<z��4o�;fY��&-���=u%�<cɶ�j��=�1�=��=�"������g�<����݅�����zC�=�<�_�
��ܘ=���<"_:�38=BF����߽�@�<7*w�|��=K��ī�=������G�V�Pٳ�I�<��<��^�;�<��1:����迻��=�=��3="d=�b�=��'<�ʱ=�^*>P��ǐ�=�B��ꂽ]�Z��P��=X8%=k�=M9�< ��<�´<d �UsL�����s�>`�Z���P}ּh2�r��<�k�K�=���-�=ƚ�h'��p��=��������s���M����S3�����=8 ʽJ>��<c�"=Y�\�꽖�n<�B�T��$��;HI���>�����&=3���T��{�!�::�
�=R�=���=�צ=�<]������=��1��Z <y�H�	吽���;��)���;x�`���=���G���E�+�;�v=<�"��(3>: ����>3N-��8�=���{�(=�����Z�~�I=r��:x;�=��L��>���X�<�����ڊ9H�W�{^���Z�<.Bн�μ��=Rŧ;8a�<��ܼ�f���07=����=�����_��5��7��<]ֽ=�:�a%W���#<�_��ѕ<�Ua�7°��(7=n:=h��񱑼�����ߌ=��=�5��-w�;~��!Fܽ����¼2B�=ָ=Gׁ=�*z���=;�=G_��=��Ygݼ�3G=i�>��M=��A�t�<��=
�`<�:�=��=��<�)<��=�H=�]�. ��?��ӫ�	K��]�'���Z�H;4���?�W0���T�?�׼�=���=��=�#Ľs3�<�ˮ��\�=-KQ��?T=/��=�I����.=�����;Z�=M��;܃4<Y�뽸_�=[��=�缽��=|�p���<��+�κٽ�:�1u=7P#=�<v��=-��H�I>��@=f�0<pf�ka9�Q'���K�=����
���ȼ=� <����~z�#��m]��e��V<���\�+;=� �$�$�>G6��:�<�w������>�Y��mT�=otY<������=i���)P�{����(�=C׭�0=>i	�F#q=5���t��=?�Լ⬺���=a���ַ�=�{�=�����XĻ�O;�jlh<��<Җs���ͽ5��;����3����ͽ`@��8 !>w�[����<�ԡ����=Læ:�R��x�<�=<|=�bQ=�� �#m��t�O<�=��%=��ʻ�����Z9o�m����	�=�Q����I=d�>��<��"���=$�ݽ�h�n�=9��=A������Խ>^W¼tGN�Y6�������>�hR=�k�=i1+>L��=MΞ<��w<֓�;���=�b�<$=W���;a�<Hy���ͼ�B<�>��&>ǅ���;���â<���]��=��������F=n>�9�=R�=�7����U���e��A���Wm�S�Sfh��h=wu��5�=�!Y=�H=�|��.$7��'�:� ��r��;�]��"]e<��<:�>D��<�W߽��h��W�%n�W�>�==���v+�=�R�f|�|���[��g==�gp<W�c=`=�<t�ս؈��q��	�?p��r08��^)��` =��=����fkȻ	�	�6�X9�ל���=K ���IH=I��=���z޽t��=��������G��v��=��=zsn<5.�<&���o2�t��=G������c�=� �r�ܼ�V�<�2��N=9����=�s#=��%<����7�$=��۽J�=%,�=4M>}w�=E�м���;>_i=�)=�7�/�2=r�C�Ou۽R��=�]=:{�=w ,=H<]1��`��=��=�t=����M:G��<��<,Z;��s��.ԁ=gq�>\Q���F���ϻ���R:�=�6�=v��O�=�g�=���;0�W=Wx�=bq1��>yGH����<�DռÏ��Y����>�v�;NҔ��L޻Ϫ�n��;'�ڽڪ��,�� >��G�0�{��y�r�Q!=O�>u�%=J�<Ǧ�� �%��=��O�;W������=h�>�+�*��<�-�=z��;|l���g\E=r�9�PX��fw�<ҫ�B�=w��e	��n,=VZ����Ͻ��.��4p�?̚�:�����=@�,�_e>uD��I�>�pG=֑���.=)���� �� ���"��?�i�����=�͔=o,8;���=y��;>�̼������7���>��f=0{Y�-ֈ<er��	��><��:��D=sJ����<��;��=���yi=�}��� >ʛ�������V;�9s����(:���="��=��=gT�;���pL�m�.>zUＮ�ٽ���=Z��=�齱({��J	��f�=�&6=��뽂��=_Ͻw��<qܽP�=�&�N�>�ͬ(=B#�<�T�<�m�;q 5=���{V=Li���y�:H�i=���<���=Y��=�LҼ�f>i6�2��=�h������
K<��0��?�=���=�� �Bj�Q���E?�<��	=ȗ�N�D�~�g=������=I<3=h���%��<��(;���=�l��?��<�sj��ޅ�%�&<L�(=���<<t�<�)�=�1���>)�>=�$��8*�<�/�=�&�=dp">{W��������:.=@��=�_ >nT���7�<R�=�cb=4,�=��R��R�=�A�e��=�ǹ��Z���ս���=���=�o=q�����=]�Ͻ�拽ZW<>�0�=y�Ľr�<ݼ^�j�M< a=Ȍ���]��Q=���^�����b&��A����c�<����v�=��?�(��;#*�����	麃c�<M�E;����=KH=(�����>s�ý����6_��f=e�7���H��5�;8^����=B�<��B=M�׺X�&��1�D��nk�;>��½q)��|K�ؑ����k;o�=4Ns��6R=����h��kO�=cŽ���� =�0�l\�=���<f]�<�E/�2�=
ե����ߺμ=����Q��5��=��W��,袽�M�=o�n=6+(���K����_v=�ͤ���'<!��]AB<��֐�O��='�
>�"=���0�=b��3=�.�=�d�{��=X2�=۹X�qo�=��)=���<�>��W=�{�^���B]W=?�h������x��j���������.<�A�<�]����=nڧ=@s�=}�(�Zp�=���;��:�� >���;���]g����ͽB/�������Z=)��=�5k;�����G;.4�}�6��:]=�Ɯ;���;�	+<�0}=c�{=��=��n=~��=4��މ�<B�=�1R=���=v��=��Ͻ� �=�l=<<��mԕ<a���E�ź�1���6=�aս�Lf=r�<�s�Z�ƽ�j,=���=OX>n����-�={�>�0=� ����=C����4�D��<��	�	��V$�=g][�A�=��<k�཰����<� >�o4_�4�G�����w�=���W{H�CC��h�<}�d��@�=80z��mn���<���?��UƑ=��ٽ��=�ī�On�"�kϴ=��׼������=(�<]�=Ŀѽ�����N�o* ��g����$>�1�@�=Ԡ�=2n�g��=Hu;hZ��6���|�=o,��C�̻�'��#k='��I:�=�r�=��E�1�;��j�b �=ȫ�8Å�=�2>�\}���<���/O�= �A���.��tr�
� =DbK=*�=2�e<Z`�=����ݽycw<�ig�	��=��<���<l����~���Y�W
>��<��C99�z�(=��ܽ?�=.�<�=�Ę����B>e�A=�������=�z�<&�;�j�=���<$����ܐ=�gh=���"��k=H]=_e>��ѽ4�����gֽ��Z=ũ�<�=��=O��=��<I�<0��=�@�=�3�=���eH=���:l��=켕@н��+���<��ؽe��Qj<g��<Y(�={�=̣Ͻ�ߡ�����E[=	�=܍��@|�=,���R;¼	�<ݭ=��`<��y<~J5>?2u=dp�=&���z�< t)�'t~���<Lw�;+^�=�"���=�޽'L����=*��C��͍�d�Ļz~=�>F=g�<������1�3u6�?�<�|˽_>�<8q���=uL�<�l=ӧ3��,0=�D3=Q|<ߟ�bvI�M�����=D}>v��=�V�=XM���
�<gs�B�>�N�<���=V�3��5�<gn�u��=��<*C�pbF�7���g`9<�=�e>�˅=�I�;�=�{���e2<{k=%���<=��<+פ<�ӷ��0�\h����p��>����*V�=�Щ=pp����M=�;H�f撼�o0�=&��/�S�JN�=�mJ=��-��<oB=��o�I�>���B~;���=�٪=�7�<ڂ=���W�;���A���8�ڼ��/>Ǟ�=��y=�
�%(
���=4�t =[0z�}����=���ܜ�=���Es=Kͼw�ҽ@��=�Y��+��=�����<~�=��{<G��{Q�=cr5��	=�m<������#=!�+=Z�=X�=I���f��=U�=!>{q�-ve;��<�(��s=4v�=O@f���b==�
	>�T�=ؠ����<{'x��r�<N�,�;f�|G�<����+�>n�o=���=!&<7����j=r˼� aļ;(�}��=DC�������o���i;�e=X��<��̽" �=@��=�=ՠ<>�s�k�o=-��<Q��=�Uü�@�<�q�<�j��lDc=���=Tf�;���=dv罚e<�])=Py>���=k�=���<���Ǉ=Bt�=0���7
�J��翼�h�t<à=z�=�{潔u���<y�f�7�!2�=M��=�?�=@=�Ѥ�U+�� <;��<��=���;�>�P<���<M�񽝜�; r��z�� J=T��:��y.9=�=��<����n1��'�=����g��{&>��:>�G���վ<���<�r��]7�#hV���=yN+>�>���=a��<샧���<h(:�>s���(=�h�9pʤ=�;>��#�	ԙ��O�I�;/Js=2.��{]��{��=�Ϛ=�C/��
���^�=۰���S������<�$g���=35=pԃ:��ƽXX�[�����ҽD8�h��=�)^��L�ol�=G��=�b';�t�<]�=zh�&�Q���5��z�=�uo��#|=Pr��	��=�й���.���x=��?����=$=�=
�<�C���X�<�)��Lk��<�hI��>��;���`T��i��ה=�R$<�>�����&�=f��={<ͽ���8X�<�N�=��=k����W��g��=ھ�=����]��
-�����6����<��e=���g��m�=1�5�=VF�;�S��"���9ļ��x;$.�=迿����<Q
����B`�<Í���氶�&j�e<T��3=�@
�__���s�H]w<$��=�I���(���v�<i��=����-�=A���Gٿ<��Ż�z�<��=Ь��U
;I�����śĽ�%�=i����=���^�?=?H
��/���=MC<���D�������y=��>G
�=�E��-����<2b���D=ۻ-�J2�=�
�߹�<"��:��ཽ}��}��I����d�;�֐=�ƥ=�� �?#k=A6��ZM��5�I���=#��(�
�ĩ�<�=|e�=�F�=��@����I>G�i��Y{��E=�����������=���3��X5̻�;>=k2=T�=hv�=��>���!�=12���:��K=�~0>�zͽl��<e�<P7��j��Ye]���1�Uxҽ*�0���̽�ɒ�إ>)Q�=$zϽ!Jt��c�OCֽ�BK=o?D>C�����<9�3=�H=�۽Y܊=� b;DB����d�xEn= \	>?8N����=P	<Վ�=�z�=�3{=0�;��;��������:W��<�I[����=&;{ =$v�=ʍ�=a��=<!�1/-=�<۞�=�}=>��ہX<���=o��ik\��*����,�O=�c�=����J������V�<��h=+�V=�M�=,ӝ<8Y�;�Z�=��> L�O	=%��:Q5h��Vr�@���c�<�>~p��I���K=�L���W=\Y]:��=��;>�̹<t^�8J=кy�ى �ݟ���������bv�S�<#C�=iM�NM�=���=�4:��=�X�=�c���[[�tM�2)x=rrֽ�W�=��X�)�<8��<�Db����=�x�q=л=�~½E���$Q=�	>�3��f�߽���;�%�x��",�vڽ�!�!�<�}�P>�g�<�^@=ǎ���t��m=Nw�=�U�;h~��m��K`��y濼�y>���I�w=Q�f�,��"CI=�͜=�қ=�D�=�@)��d>��M��=�޳�S��< �=�~���چ�L��O�ԽCUν�CٽR�R�h�Ǽ+�����=������n������j=웆=���=�_=��㼺�z��$�|=$j �G��=C� =�^�+�½�;6=��K�OE���冽>�<&b-���;�G��ϓ�<���ֽ_��4g�#���a˼1(�=��<�-<�@��V=��n�b�ƽ,]�=��򸱟�<E9�={��MR<�(7�T>��ږ�=\4�4�><��o=424�T�˼��><�M=kTH=�	�;M[�� ��=[��=��#<�a�=Bn�<7�=q����=�$�=�9���jټd��;�L�Bz�yw��+���<u�=��L�¿o=6�߽���;,�B;C���e���=��l=����#r���<�>��0=Hg�=+!1;�y=ZC����2=n�4��.�=���=�V��DŽ�`�<H��\#�<�S���Ż.�>�V�<�=���<�=����E��}=;�ƻ�G�=d�<���<A�>)I;4�����/!�=�*'���=��=W�0�M=n�ɻ��<`7���7�일Y�ݼ�"=�z=ix�=3�=�>=N�p;�S!>���=�l";���<�(>#�"�C�c=h	����<#è<=x]�L��=S �<���=��X�֏1=���=�0����]=��:)��=g$>��a=�i\��pɼ��;�%��ͮ��ký1����Na<�<�.
>�Ð������Ѽ9���l�=��{=�,��@
9�������\�H:���D�<�H�h@����=SB�t�z<O+��/���ۡ�iA�=�J���;K��2�����!3�=֚=Ri��ҿ=S��=��<�a�=а���Z7^=T`�;*=�==Y���-f�y�;��нt���O!�|�7� >,=�o��B>�<�<��ν������;�ɻ�X�=_/����F��a�=͹��&*>�S�� +"�������=�Ǽ�b<���ϼ�4���E����=��뻨�{�J>;��ܭ=@��=��=�i>�a"�����<��;0������ڛ=�7!��ݼ��ֽe�<��ͼ�1��q��=\�u;�J�=m�;cٽ��=���<)$�=�1���ݠ=�Y=�P0�*��n��<�<�'A��Ѡ����<��'��=B)�<��=u(�=:`+=�o1<ˮb�H�=��Y��?�=cR�=#��<tٙ��r�����=ew	>�림/|�=4=�=�*ܽ��=�N۽΀K=�@<�~����=����>��=���=�۽$��������=��2�c^P��+<�%=�h">(���:��ҹ�:O�5=cu��0�=g}<�G�=w�=C�<��<��=�L�= �=>�t>!e�Fio=�q�<L��W� R=پ�	q���E >�+��(ճ=�M=w��'�i=4/��^*>��=j[�=Gp��e�<É������Q�"=�C(��_�=�U<�{n=��=#�B���6<͊(��5>�o="�H�����t;; �/ҳ��ZU<퐼�d
=k���{�=�ٽ��2wٽ��	=����r���L�p:�t6C=c"���%�c�ѽoR;�Ĺ=�z=����;=����2�iD=~ѐ�l�����&�=�.~=
W��
>��<w�=�o8��و���E�=E��=uo<�����>��˻�ۀ���E;9�C�%�������'>��4=t@ǽO��X��=�ے=��Ľ"7��S���9����,=���<5v�=�t꼛	���,����=��	>��='��=̉�<p`��`�Ǽ�w�=H���!U�O�;8丽��Ͻw�ż%	>x^̼Mw�96����=t�����G*e�R�Z��������K�=|<D��<�t���E=W����=�M�������)�=��#��A7=4��;0!+=զd���<l�`�ݻ*�X=o�K=<\���=#��8Oμ��C=i1"��=��ԼL�/�����(}m�
|<�b�=o'j�x�]�Ѭ���W���'j�G&ڼ�I��#߈<3�<s�`�U��=T>�=b�>��"��j=ȧ��+z��w�"<l�F=�L`=������xD�r�g�8r��O��<|�K=��.=aD+����9�:�2!�j�=^T�Ҁ�;�ч=�$�<������:�!=��{=�n��(d��i��u#&�vk�<h0!�]���Һ<,KM=��=�0D���=�I��w��<��V=B����0�=a]�����o$=o���N��{YA�s���F�=���s��{RʽK�=�<ɽ�R��-:)<`�>$��=&8C����L=<��a�c=�Yc<�m�����=C�鼝�i<���<&j���K=�	�|	�I���b�=.P&�ѿZ�x�<lT�=�����Q1��$�=� �=��>3w�<X$>��=g<>��<�*�<L6��P ����e�Ф�a��=���;x>��x�À>v>�p�����1���={a����=k��<wA�=҇{�G�=�a���e\���$>�@�<�L=3O����w=8Sg��n3=�N>Q�;����q�׼w����z�^ͽ�����H=�?�
�����~=�Њ�,����l�<#�����~�̽v$i=���=��!��^���mM��>�ik=���=$��=�;;�4�I҄<�񼋩��6�=��;�?>��>P �=0:>�{]=
F�=��=�G�=ס�<?ང��=t<�G8<��= ?Q�����q=A�|=�BE�1K��۴��#���=��=3���5^=˖�<�L���j�j��3&w���/����=��#=٠�=��!<WI�=t�����ʼ
|��pڽ���;<�¼�`l<6Y=	��;2���D�E��b�����<˘�=`��=IO�<Vܾ=!ͬ�%�L�_x=�zݼ���xY�<�e�=,�<�F�Ί3=iY�6'�;m[=+{��F��>�.�=T5=y�=�I��&7=�6+���,<$f���T��K��=����&/=����Xڪ�v@P<5�<��D=�N��'�=�P�(s.=���=F��rԴ= ����d��U\��M�U6@�����*��������ܼ��=_ȼ᠐=���n6�=d���{ <���<�{�=H!�|�`=�� ����=:�b��Tp=�$=�p�=[��<R0����=AS����c=�c��F(=fS&>_ď=�{��P���4J<`?�=����ń>�V��������?C����f��Q����<�Xo�e"�;&t<` ��V'�D����ݽ�}X�nl>��ּ�*;�Kn=$d��f=���=ϝ,����6�9��?=}��<�TJ���=4k=�ڽ���=]���?=�4=��=^���4=']��<JA=�l�=���=1�=~��=��+>pȑ:"�j=���=�����=�p�=�L�1}=��C�2n>~J=�H�=�`e�:�	�`�Ƽ\�0=�o'="�
>��Լ?�=�t"�q���+��5�;�D��*�����j��#���y�<1��⦽�n�1�򼉲�=�U=NWz����=�t�<P������<�$/���F=�;�S���ӈ��n����<��?=��u��=�5=��\�l<5+�=Ŷ$=�R߽�+>�=[t�����޽">`^�<��B�,>� =A��=j�=l�����<3���&��b���TSp=(֫=Ȉ�<�ä��˚�ՄW:���g���}�<��A���˽"����>�ҭ=�n&>k���4�˽�T��R�=���<�S�={�=�E�<��=���m*h��I=>]"��4O�j�=�<�����=-�u=hC����=rCT=%E-=F5���=>�-�#o�<�hսf�
�`W����<�3û��;��X=��Y�9)ǽ�ߏ��C<���<���=3.���Z=�;�I�*�j��=��=��=m���f���8%=p>�*=Œ��o�U���8�*$3>8y�<�GĻF׼�C>�	���p��ڵ�=j��;���=��!��₼�ؗ=�%=g��@�=w>E0'=��=�P�;x�T�M�
�w�=C���Xk�Xͫ:���=Y�:=�Ə�pwT=�v�=k��?�>6��=�Ƞ���l<�7���7��)��z���M��=E`=�6�<��`=	�����=�k�=�:<9����z�=���׆��S���μ��x</ڽ�K��@ݼ��������J�3�L�2�
>D6ٻ(�$���K�;�q�=��>�j�xѵ��ѭ=H��k�6;��ǻyg�d
<��9������=�
�=/r�;��,�>�%�Oؔ=�<�l��B����T=յ(=^�<٫�=��=	��='A&=���<mwD=.��=�ڽ���<4;��H9��mv�����v6.=��>R�=h���3���-~]�A�V���=�H��F��<:�����o=��=+N�=!�j�ǆ����������=�\�<��x=󲉽ƿ3��㩽7ns��Ғ�ܩջl'q=���>��=�������Fw�=D'=VWͻp��=s�ԽH�^=ng�<c �=Ns"���a=�3�=O/ϼ��q[��ڼ���=��<�_�=ڏ�;��]�޹=���ý�I���zE=�	��G$=7��=G<�<��l=��u�Jv��x��=��9;59=߰��h�=Y� �J+�=�]=�����U�=���g;��r���KGi<|/=G�%�7:��QG=���=TCV<��y�}w��5�z�x�h=3���A#=���Bz{�0�c<yhp�bo����Y�)g������QF�6v<�k⽥Y��h��<d&ͽ$��=��̽��x=�˔=�|C=�I< T=w��=uW�<��<�B=-�=^&-�V81>��=�r�=���<�s�;�����
=4:>�(t=�?
:̛�<�o0>�$���`��j�=i��=��5���Ͻ^ C���6����=�l-��U;���<��B;x�/>�'=F�T=� ;-V��aD�<�	�=�����Az��5�<PF=�8=����41>��<��<��P�>����<��<����>*-�<��=����3��P�f�
:���o�;;�e�M�Y=����i�<�l�=>�=��K��F>ّ�=�����~r�+�)=\ �=�y�=�᯼�J�3H�=>�;�>I���nC<I �=��L�4�I<��=[l��U4�?z�[�ݽ��D>��t=�O>��r.�=��<�gs��o�=|��<��d�ֽ��l=GGM�#��=�`�=��C���$�E��=Elͽ��=��>��ӽ;"��}O=����>��<kG'=��=M�����=+�[� ��5��T$<Հ齔ؖ;��=H=5m��,���;�2���n�`�H��z���<��\�s�����_~���8���h�<�E�<��6=�u��ŷ<�w�<l޻�q<��>=�	8����=O����\�<&뎽��J�hy�=��=z��ę�<8(e=�j��r�3= {�=<T�Z)����=��^<�f��<�<�N;�1�d��<e�s��s3=�a <�>���=T�=��E��<��R�=3�=�M_<��s�O�<F#��6z���Z=��S���<	��=\��;�����w�=�*�<�
>�I=�,��v>`=����=�#��l_�=��<�e�=��u�w��<�Ʉ=��\=$��=�������=RyB=2F�= #S<'ͽ��=U��<[�X=���;P>hg0>����\����=�
=�T���Փ� �u��Z==-���
>~��=Ԩi=2�=#��ᯂ<ژ�=�
=!4U�`��Ѳg<�b�3����=�fH=ɀ�=r<�=�Ǹ�l?��1w�nؗ��¶=���=ǣ=�޽ ]=��?=<�4��$>0q>��%��W��3�=n�,�>�=4Ԭ=������=��=צ�8��=�u����f�}��:M���2�<Ѽ=Sx<�̚=�0���^=d{��5�<�����j=�𔼯��=-<���wm��#�6R3�h��=靬<=4�x����2U����=#]���n=f��<�4P<�����	�=� ���ݩ=��ȼ҃����;��ͽPӊ���=�н=S	l�ǒ½9>0�Dk]��u�wA=u���' ��=�&�=�VY=�`�=bB.�m��<�l��ya�\������=�%�<!_�<"4;=�.=������ټu=�uk=z�D�����&j<��>������dŽ[*������;�������F��=��V=T�u=>�
�U����"|=���<�ټ���;�~�=ޣ�=
:r0�;�1�����=`o��v��=�}����>=.��=��=��;�%=i,�<�ef��q��YE<�%��=˓�=Uh=�|�l���ƊX=Gսy蹽��K=������=��> ��j<�;�f1=hM=�?�<�o>��q<�����S�2����=גB������C�p
q=��ս<�]=o�>7�>8�>���	�@�9y=�.�^6���=	�g<*o��{�=t�(����O%����=Ǚ<2��A5���+:�Q���z�=%�g=�����p�n9�|Q���!�<�J=��2���������Z��j�ܼ0��u{���%���aR='�����={�=��ѽ2�3uq;y�ƽ٢C�v�v=j�ǽp�̽��=���=�9�<��P������=��
=��˽��<���3���䲽�!��s׿��>Q7	=��;>��<\��=�̞����x��;�+A����=�п=urn��i��\�d�2B��/��<����p >��ػ��.���<�g<��I�)=)=<tS��^=\M;�=ǽ�߃=hj�=3N��"�=��=!���E��J�<([='��9�@h=�7ۼ����/Y=�>z���=ڣ=pq��3��t���M�� =(=��=޴�<$�u<ؽF(h������M��25��3�<�Y��ri#����Q>6/J����2	�1
ƽ��=��D_���ҽ���=s˱�Z�E!�=1b��:�<酨�:�>�U��E4'�6�	=ԑؽ��l��L �A.c=Z犽?Q�=<{��aB���%�=��<`�K�!��<5�=]��<��<�I�vg���.�<�:�=�(��F�d<���⪔�����wG��'�`8F�a��l�=�r��A��yD=��=�����c�=�G*>�k���M=%�+���ڽ����*����<�\`<h1����R=?%׽7���l����g�r5=��ͽ(�<�w���^?��o�����;G�����=�q�<��>C��Ŕ<���,+��zz����� =5_��oѽ^��;|��=���p����<A�T=iA*=�^�K(=��-���
�;��=��=���v
�O��`��r
��;���<|\R=s[ҽ��<e�r��x2<�6������f����Z�rd�&͒����hƇ���n;Ƅ�<��|���o<�����['=
e=N� � �ὓj8=�ӽ�Ž�ֽ8ׅ=G^�������;E�J=j�=���L�>lN���V=�I=���t��˒��ѝ�V	��=�ռ��=�)����<\���>�̫<x��=���&>/�;#7���ݽ��D<$=2X=���ı=� r=`���3=L���p��;���@�׹r���O��Z=�
��l
�=v >�ѻ=?�R��2�<	�����="=�Gg=wly�1��=ο�;�Z���q�=�on�aM���=;���5�=���=,Xr<3_;��Td�)%�5�7㽏��t<�=�R�=�o�9`�&;�	=��Ҩ;�ӣ����<$�>!�p=�>��b�>��=�#;��\��=F~�=fѻ�H�;C^���u�=�p=.=�=��9=5l?��޻\+��R)+��K>��=<w=Y ?=S��<�����2<(N�����<�⺽K���?�=ey=\��<�^O=��#=GA�=�=���><�=H�a��G>+���U�=J�=b�3=�#E>�&�We���as>X�<�'��Uݽ�V��ᬽ@z�;��$�	���pq�=��ҽ*=5><�X�<�^��qz���>E!�=�S�Q[�sW�<*G=��<�컼!��@E�}�=���=k�<�3�=�9<�ߖ={�
�i� �A�V�(��<f�=����߻iq�̈́=YL�=�F0=}�>��{?�=?zu��#�����=�5�_�a���� �(~=
��{�*=�ܽ���93�
4�Ac�����%n�<���<Ք>�U�V�,<1J�=\�?<�|ֽܳ���=4�ƽ���=�O���3B=�J�Ǵ%��W���������L�����=�N���漰�5�����%*��,��=B��K]� '��.���'���&���=E(b=�9?=a�7/����=1Ӻ=���=;�<W1=-������=�N׽U�S ���8�=�ݼq8ɽŰ=�&{��~�<Lz���!��V��=�|����<}E�<#~=I�����=�1�=�<��|w=��˼�6�<OQ��~�<�-�'y�j�*>Q?\�<��=&�?�:�.��l=��<Ϧ=��0��p=X�<�{M���ɻ�p�Z:];�l�=��<��M=rʍ;�q���o�d�=��$���z��Q|=�Q��Y޽��=�	=N�=5��=in<$#�=�b�=�+�=�۩�<� ;����2��=�|=�Š�I�?<��=4�z=���^
�=�˽aC�= 
^��W=�1 ��
V�7Ȼ=��>}�G�7 5�;-=��;=�qC���<<��=�n���޼ �V�4r=ï>�x���#>ldW=���=1i��f��IPY��}ں�=�xO��E���ܼ7������={�=��̉E<f���.-�]ȼ�;��`���<���;>>�.�<��+=ң��W=<�[�qȴ��~=q����6=���=^�	>e�	�
�T=rk=�7x=��g�>lG<m��=3�ܽם��)��Q	,>���:T��<����c�=�ױ=�C���=Z=E��=�X�<LΥ����<��=�#���>;��c=ϰ�=�-P��|$=H�=#�&>f������<��
�/;?�>�����=<G��<��U=�L�=�)=ǖ���#=`T�=�	�⽢����=�����=�=�]=�s����&�g�=،�\^)�a�:���<7��=p#�(� �����=m���?�ŀ��iP���<?wC=j�f=��C=t�2�0��=Hz�=1�Ľ��(������K�.��<l�ռ-�J<6�-����_0<!=e�He�=;���»*�x�G=���1��x����#=JO��Ec���L���|���m׽&WB�a���t��
��lτ<�/��s�\���8���C ���{=�w���S�������E#<p6�=�k�2�X<�=>�=������#�
=��J=��:N<*��=2:�<̀<��=����r���w=v�Y2������>��>f��������,=��~=��=��S=�L}<:2�=���=x�0=���<W�R5�m�N��,������!=��3<��=��=�A�=�_�<�t}=�sr=��8�uv�=�x9�� >�3��W*4=C��=EW��� {:�(7<AC�=�>'˻<.�M=I��e��\_�=�A�=8e(�/]�<��ڼb��=p�=���<ؚ�=ڑ	���e��Ԑ��Fƽ-�� �
<g�=m:�=ӺY=9�=�0�Nz>�í�dט�V�8>����?Ļ/��;ʌ6�)���ą�����Q�=BǸ<�%�-b�='�ýq/&��F>�O$�X�H=�pѼ�x���=�D=�᩽;8����<C=��лp�=�!=(�%�L�нk1m;p�=�=�B=��5ؽ���=���2�d���=�
ӽX� ���P�F�<x�=x���ݙ�v���WƼ�5W���>=����(�=��<�I�=�R�=U�<�_½�q� U=u�=s�$=c����<��W�)����@=FtM�\5�<@�>�M�=X`o=�����>A	+<�h��CV��c1���t<Pٽ�fF=/ʼ�9�:���=����~c��T��=x���hU=�J߼�g�=�)��hs�Jýx�q=Vc�ٔ<�ν�0�=���;���=-��=`�N=U�p��a`q=r���<�8������=�c��%�b��]V�;)��#�.�=\�s=\�ս��=�e����>�k<�e��X���&�*��=f��Ӗ>�����A�/=��4�=��]�X̻��U<L�.<@V(8���<p�=W{�<q��<�X�=痹<�M���;'���=g��"0=�=�	ɼ�c_=�=E�z�� ����<�ڌ�}eM�}�L�ҽ���FνL �<�_�<�
>7<�=e��=2��?6	�	9>�޼�59D����=&��=Я�=X�<�(�=�?�<c'�< �=BĀ<�
�=�!Լ�=Jߑ=�ْ=���<��<�03��a��X:�<>۽K��=Ͱ��� >�q�����)���h�2>�f���K���<_)�=(�;3Ж=耼��
�a�:X~��n�.��=�J>�������aǽ��=��d<\V��ş<pY=�J=��.=����Ǽ!=�(���a=��=o'���>��̽؋��j��<���;���=��G=��o= 0��u�=q��(Z���?�����n;�$�_�k����<�>I���݁������G�=� &<�1L=HN��I>�<������.>!�Q<�����v>�@�8P���[m��5����<�-����eO�ep�:~Ow���̼/."=Q��=��Q�G��h�K=���� �(��=�R��:��<tmk=�ɉ��6>�ួ��I=h�<���=㧍��������WK:9nԽ-�O��N�����o8� 9J�9��\:��ѼC��>�c��m�=�2=�����P8�B�L����;�]���;��E���x�#Ə��=��p�@��=Ӡ��}՞�PWڸ~ޫ��<�ᵺ]=D�=ǂ��<�=8��d�<��=�~ټ�ݛ=V�#����=��<ڙ�=��=��E;޳ ��H��������M����=RŊ<�1o��^�=�1ν�Y'�U�+=��<c5<�P��4���֥=Eb>EǮ=[�=�p�<��<<ix��iX���0=\��=��他9�b�Q�2��g2��O���[=W?��^�ѽٌ̻��H�{��=���Nw=����zZ�HG�;c�s�W=�=`���P��b��=�G�<�,�+�E�h�~���=hJ��%��Y����R��d=1�
0ļ[h�=2=�É<:�(�KY=��<�;]U|���s���=L��= ӕ����;^Ś=�����𿼴��������`�� >���؞=.��;�&��ǵ�i�)��9��->�`J��R׺{o:>�{9�B�L���=aXS��������1=�v�=���=�i5���n�K;0D������®��娼�ׁ=��)<w��=m��<�W��
��<#��'M>l�ۼH:>���=L��<q�<��=H���8R�{gL����<�uj��}��l���.ѽC��=�/���`=_���p{ܼ����Uw�[̼+HI=���>nU"<��u�H�L=T����C<��;(����������=fm���
x=�\Ͻ�>H�n����:3��v�=�I>��U=B;�=0�%�M=u�۽F =-�n=���2$ ��CV�>���w4v=���=�^��ѽ	��<���e>=�+=:r]��ͽ�o�=o�e=TT���zT�1<�=�C6=EN,=�:-=ߑ�=���H��mm�<>p��G����RG<G�=F�<�;�=q��<j�U<ງ�FOy<�z= 	���h��4��<�^\=\�?�c�>��}���E=;Ʌ������='�=J����n���*��N����<�<�$��Q�=���=-�>�p�t_����@����뼠�����&g�=�K<�H+�����Tǽ�r�=f���q><���_��<Æ3=i{8����=ǧ���y�=u�<$�s=�P�&�廭��=��=t��<8���?��.�=�I��9߽��v=�̽諼�><�a�<o�ǽ���7�=Ed)��R	���ʼ���<��W�9L>`p=@Ml<�C�=�?<���./=�	�=��= ⽥�c=sA_=屏=�%1�������z���0=���ɞ�q��<s,�;�� >�P��D�^=������N5m��	>�qI=�A�>�)=�>�f�=i�%���C����<���=�ef�B�I���>8�������ʳ�ڸ<HX��J'�=/W"=�"�<dU�=�1�<.6��֕�=(1j���=E�n��J>=#|%>k�<���< �n=�ļa)��GM=�����'��=�A=�����A��=��<�������=�u]=$�n�40�<eV=�|˼���!�{����:�RMD=V�>'�=������&��������J��Nm<<,�r��I:=���r�,��˽�I�;�:����=P��M�����=c�=��<;��<I�;=H�꼟4.=�(�=a��=)����;��=*{�=|r�=��Խ"���D�ǽ�a<=��N�@ㆽ����9��<3���$;D�fx�;�x��D�¼B�gg*=�獺,G_��{=:	�����<{�<|�н��%�W��pU�9�5���Kl<�⿽%���º<��A=�����b=>P��xi�=�Խ�J��<Z�����Ϳ�<p�=��;<��'ҽ��;���,=)-=App�H�X=}�:=�ݼ��=v<�=j�=QQ$=�-伊tG���}�<���=>��=�@�=�0s���A��ؽDl>k�G��.����K�=�b�=B*�uNݼp�y<𿐽��g��{j=��V����8u�W���k�=�u>�\=$�ֽ��]�=;�J��<� �ҵ=69��x;���<�����z<#=i�=Zx�;9:>d$,>ބ�=}��<�a�Z~O���;��ļZa�=�฽&�5� /�;�뱽�$
��G=Fiy�*M��Г=	q2=!x@��y�<ս�=�d=
(���=�o�=��<�7=�!�����R\߽�?�=�)�= �0�0�_=k�=��;<R�<-�(�1�<'��<�V7�N�6>O�=,(�=�v��)�W����S=�r�=F���xr���<d���=�<<�����,=�Ӊ�:����m5�gz��K;��>�/b�߃=�T�<Z��=���;��=�Vx�y�=����=��>�d޽H�J;==[>�>��>,��<4��=�X0��x��yL=#�=>�~=�b�=���=��>Pآ<Gي=-�<��=<=T���ү��vҽv�={�=��<��=���u�=W�5��59<��W��[���s��=8S�=u���������b�E��@P�� �=�5�;� l=b�>1��=:@Y; �Y=[R=<� J�C�>�#"=��=l�;	 �=nl�:�E>�4;��l<�ڻ�@b�G�
�d�#��=~P�����=q-��r<��<e/h�𰬽���� >(8�v�=��
=#̫=�JA��5曽!��=�H<��<�t<|D>E��<x�K;��H�Ɲ�雇�ΰG�2�7;�i���R�l.�=/B�=��M=�K1>���<b��<���=�h��E�e=F�*=ڡֽm5�=2��<��P=H�<M�_��oN��7O=��=wk=<:�>�K���D�<���<�N�3�V�೽�׽G��>jZ�j-��{p�����<�z�=<];�dL���<��J=3�1=L�L<٥�=bm >3��;����\���c�Gb='�ü�z>d��<u:=����1k<�:<\ƽ�X��:���S¼&=��=9��=�I��^�h]�;oH>�VϽ��=����<�N�<%���\�=ܧ=$������:�c%���#ʽ��8���[=g���ޭ=?B�=��N����=E�=[��<�]>&2�=m=�7��"��'9�<(=��>=N��=H�=�E�=�`$=3�=���=)W<�臼��4<�r��e��<{�W����<
!�<(�=�~��j�=(���=A�;��,>����'=E�>nׯ<�z��{=�F�=Ŧ9=G�=1��=����p=��;&>A=���=�� �9dc��=�/w=�z�=g�=.�� �=+�L�b��$��.0�<ƞ���<�_$�v�'<j/��k�;3���ZO=�A@���	����p༙ƅ=j�ҽ��ȼ�%�*0�<��0=�Ǯ<��{=�<��h���N=~�����J
1=�*B;�V�=rc������>�Ɋ���=[�=4�)=B>�lJ�*zS=m�<�� <����5= !��0���K=iy=u׽��S=R�>��;�!s�q4Z=��>��ҽ��=+?�LV=j�->�/�=M{i=/�E=/���y�=�)ؼ��W���r�ɮ̼�$�<ߋF��a�=ȉ	=PL�=7�=(e%<��9�}7<�d/�u���`e��߈=��߼��=nN��R�;�4�Q~w�A�-���<�8�=d���X��<�=?���4��=�M�=!򼰜�����nN<.5Ľ�U)=ۄ���Z��l��p�F�w�޽�H>��)>]�<�מ=����=rT��>��<���<��=zIݺ��>X����C=d����H=ܽ>I��?�4�
u�=��8=��!>�G��o��"������	Ƭ��_�=Ih<II{����=�P=vHN=�!<+սt���Y[=�>3-�;��#��8��R>�K=���=MT�=uX���J$<�9����;���(C��
��������[=��7=��=�Ƴ���=N�<�r�<�ϭ= fn��#=�u＇7x=E��<�x�;���5��<�[]���=
��2)='��=��2���j��E��!�=�������~�=��=/�d�! �O�/�07�=v��=��=�=>`��6˽�=*�<�U������E)$��bE=�����=hJ����=��Ͻz�����~�w總�]�.��<�#����@�<�Q-�LM$>vX:W�>l������=%�!�
�< (��T��gjw������:�<�|�=,%��?��=᭠�չ=o�:����X�=�kѽF8<>׆4=�P=���=9�v���="��=`���pu�=9�_=SR�L������<�,>�9�=�����R�X���:�o�q��$=-�J�e�nހ<C����L�=*��ꏻ�.2=��ʼ�z �����N�=��n���]{����T�ӺW)�=��%��<L�K=�Zr��:��x>v"=�V����y&�=�o�sK=��=6�/>퍪=�?�=
��=����u�:�*<Z�#�R����3���=#��aH����
�=}�<���p�!=��=E�Ѽ�E˽����g�W����=���=I��=ԁǼB�a=�w�=�a�<�5�v�+�sdl�i�=�ck<�p.�����^%=ɻ�=(���ǐ���>�''�)��<�f�������J��M+��T=���=^%(=1,=�o��k;=Q���7�Tb�<XT����g<o��t.���΍=YAI=���=�⥼ѳ��hk=������C��?>�g��*Y�<��ƽ������>p'�A�0>s�=O		=�Ś���=������O<5���2/���B=�L��'�.r=���<��&=�K/>Jwm���V<*� ���L�j��=�N�=Q�ѽ��=#J-=�x=A�/=@��<9�����<�z����<������=7^G=�㶽`�">˖=D��}���ʟ��t�=�S��,�i=�r���< ��,��s=�Žzj=|.�=�Z㽅��`O½��>�R����׽���B�<Ih�=�`d����=2DM<]{q�LNL��
�=7B�=�����'F<:p��ݺx� =H���A���(��bͼ��սs���'��n�����Z�S��"�<%�=�����=23���������󽭩�=j�=Ԛ\;{��Q�v<`��=�\����<,�'=Y�!�6�����>1u���ս��4=��=�~<��@�	�X�11\=~=�\绦L���&P��:�:��->Gc>ӓm</s��8��EH]=�y=ྻ�S<U�;d��rK����2=�0޼���=�B�=3��x́����Rϛ<��=�e���(�=3qS=�ѽ�>����%�	>U�=��=����a�=B㔽��=�ʪ�����D��A�Q�F�t�m�=]��<ʹ�=�Q�<�3	��I=[��<�g<��ͽ5�{<���=v$��Ln�=���p�e='XW=>}��Ɖ�ƥ=6
Q�QBȽ׷�z?=�MM=8��=�L��a_�9N�<Xf��\ŭ�Mri����=߃׼�߽)G���V�=�>=5�==�B^��C.=�S�����t�=\3�h !<xj��(
>&q�z|����$�e�Z���<M���=��P�G=Ui�<M�=[N>�"��g��=��Ԃ��;�=��=�'{=�E�=qzU=]���v��e�6" �)��=Ϣ�<J�0<ct��p@;2y�=�a=��=S厽w�.=�X�=j =)�Q>�x���@p=T~�.!��Fz<�+t���G��fZ=�w��f|b<�7��<¼s��=��j;O�h=��`�3��<v@B=��n=f�=Q��g{�<3C1>mU��+��Ds�J�O=�P�<x�qX\�ۦ�=!��=z��=�<:����q�=��X=���"1S=���u�� *=6=�{v���=��u����A?�=�ح=u��~�<ܾ�8e�=Ms�;�Rk=�<��#=���D���F
��?��Y�<�	=.ʛ�x��<0�6��>nǽ5g��׎D<�1>#U	�:�����޻:��=d�1q��u��=y!h�(=V9)��r��Vd)��q�����I=i�=��<���=J~�=���T��/�μ��M<u�=�ս���<��='@@:yݼ=Rb��ͩ����$n�����K>��=�Z�=|Q�=I\��0�ί2�JQ�=��߼��[����t��&*�.�;��p���)=�i=��ۻ�y�<���=��|=�a;T�
=c��[P�<�)J=�)Z=���=��=PA�f7$�����Ga=Zv=9�=a!Ѽ��=�p|��h >�1�;�֡=,���M��=]0���)�=ދ2�9�����B<�<��L���ͦ=3i!��=y-��gS����ѽ�oX��n�=:�̓g=�i�Ĳ�=z�c=U�߻Ņ=ծ =XC9��;~޽��=A!d���9��<�&H�}�>x7�=��a<����4�E�<��ҼW�<�ۺ=d��=zg=���=� =<
�=�0<���B?i=j; >�H̼e��<}�=)��M��=鏽?�=�7Z=A �=WU�=�)=`i�=bS�=��=xBS=Jt�=��ռ���K�/��k�4�=&@0=�O�BKN=�=l�= J�<��=�_�=|����,��&�|<hP<���<�{=�����h�g�>;3���)���7zW��B����<��>׵(=�d$���ļ�$T=�=?���S$�2�<ȋ
=b�������ꑥ�uU>��3=�Q����7Ó=]��P�<q�����=Xc>=�= �<�=>���g֒;	Ɨ=m3���
=��;�$�=�4��Լ*�H<��{�v�ʽ��>ì�=�n`��$Ѽ;�=��;�^:�={������8�J꡽os3=Iإ<n�0>t�>��O���� ����=CXٽ���=3�=��,�N�����>��)����;�/��<�Iʺ8H���z�<v�=@���$ �ʎ�<I/�=׶Z���G�[�k���=uw�=�$>��_�<i\���6�=_�b��Vʽ�	O�b�w<�fν��<�_~/=y.�H.�����`^ż<��99�/�ǽ���=0�==���=@�!���k���UJ���*=N�*�Ɗ
>v��N��d%"<�J!=��9v(�=�=�f����<$���
4��>J;qȅq�Rq�K KzKz�q�KzK�q̉h)Rq�tq�Rqψh)RqЇq�Rq�h7h)h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222174816qX   cpuqKzNtqQ.�]q X   94889222174816qa.z       "[�.�=Qt���_���܇=�����a=vr���������ư�==��S{F=l,ٽ{�=l��<q?9�\���
�=�B�<� ӺN�����(gb�E֐�wнŪ���<-vk�i =h�-=Ԡ���;l�c<h
<�_�<f^=��+=xwݼX l=@������9=u�f=q�C���=�T�=��&>�L`��͕���B��_>�|ûb�>�=�Mܽzɰ=J�<�����\��=�f�q*`=4@����x=�nN���ۼ0ȕ==;=����r<���8G=<��<���=bl��-���=nI1;k߆=�L���=Q�m�fN�=KX=�Ϣ���=��齢W���_�=��s=f�_�����4;*}]=���<�V�:Ӻ�=5��}^˼xj½�'=���;�ǿ����=�����<F�Z=�fy���=�6=-K�Z=��=��5=a0���н�-d�"_=�7=qӅq�Rq�K Kz�q�K�q׉h)Rq�tq�Rqڈh)Rqۇq�Rq�uh	h)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hJ�hKhVhLhVubX   1q�hYX   2q�hf)�q�}q�(hhhh)Rq�h	h)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hh)Rq�hJ�hqhxhd�ubX   3q�hz)�q�}q�(hhhh)Rq�(h(h)h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222254928qX   cpuqKzNtqQ.�]q X   94889222254928qa.z       ��?��?Ȉ�?!N�?+��?ā?B��?�h�?Ao?��?Fh?τ?Cׁ?D�?\m?�?Rb�?��v?C`�?r�u?�r�?9R�?/��?vLt?g�?I�?��z?{�n? �l?���?��s?��?#�u?��?��f?�&f?v?��?��g?�u?�W�?췆?s�q?!ǂ?�=�?��?J%q?8�|?+څ?|�?�q?�m?��e?�l?�Yr?��z?S�?�h�?��?�Kt?uy?��?�U�?�Mh?%��?}�p?�B�?K�m?V�?�{?�_v?qrs?�ه?>j?Q�w?P�?�\?��u?
��?
��?��?��e?@|�?_�j?	m~?�~?Tzo?��?��n?�ӈ?]�}?�t?��?ks?���?�I�?���?F�m?��?�y?@�?�.�?'�?$ w?�^�?�Fp?�8�?�=v?�u?��r?��u?$�x?�E�?��w?$}g?~�n?K)m?���?�J}?+O�?��?�kw?q��q�Rq�K Kz�q�K�q��h)Rq�tq�Rq��h)Rq��q�Rq�h7h)h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222255776qX   cpuqKzNtqQ.�]q X   94889222255776qa.z       ���)����=��l�1�m��m�=3޲����������=[��=Qw�(=���ͯ=���q>	��=Z�<���=�`����0>*+�=63ؽ����sS�<�p�o>Pe��d�̙ѽ>.	��x�����Fg>�=�=���;L>�����,�x��=�ӽSB˽&7�����:mM<�B���z��?F���Ph=��=1�>�����=k��=�Q�:��=��=���=��k��/>��=I>��=�#�=�f ��2==�����u=�W��u= �`k�;㢽t>>1�;Z��=um�=����)q=M��]�&>���=`i�������L�=5�A��j�I���8.>�:�=���=K͞�)�B�:�=��=�2>T8E<��ؽ)���������=��p����=F������=}��
;���=5��=��g=(z`����=ۣ�����=z����5���G����=r.=���r   �r  Rr  K Kz�r  K�r  �h)Rr  tr  Rr  �h)Rr  �r	  Rr
  uh	h)Rr  (h�h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222256624qX   cpuqKzNtqQ.�]q X   94889222256624qa.z       #��>|��> ��>7��>(��>�k�>�|?�7�>�a?Å�>;?Ц�>��> \?!�>��>Z��>VK�>�?oI?-��>�s�>��?ն�>rY�>͞�>��>$/�>�>n��> ��>���>�V�>��?���>���>�x?	��>"�>��?VM�>�f�>[?�$?�?��>?�4?��>.?�>�R�>�?,(?�zJ?P��>�X�>�:�>[��>�U�>�Ǽ>�h�>&��>�?��?8h�>Ȃ? ��>,��>?(,�>�S�>���>]�>'�>B|�>.?���>&_�>t��>x�>޲?Ɩ�>���>��>�\?�2�>�^�>~?6l�>~'�>��>�&?��?���>\��>'��>��
?�)�>'#?��?��>���>�>��>���>���>��>z>�>�Ư>B?a��>���>�W?6A?-^�>^��>U��>��>C �>b�>O$�>��>r  �r  Rr  K Kz�r  K�r  �h)Rr  tr  Rr  h�h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222349856qX   cpuqKzNtqQ.�]q X   94889222349856qa.z       )��>LM?���>�l?�a�>%�>�5Z?eX?$?p$?Et�>)��>m˲>0��?y��>4` ?��?e�?�$?�L?�W ?Z��>@��?KQ�>��4?�?>�8?��E>.\?��?�m?F?'��>��?���>)�?`�?�	�>7��>|��>iO?��#?e�,?E^:?��%?V�?�B;?�\'?f�?�e�>�y�>��?�D�>N�?)�>��?�a0?,&?�
?B:�>��&?@��>�S
?��[?�
?���>Ts<?"��>���>�Ɏ>�5�>�?#7�>v�>�Ѹ>0aW?*�>-��>���>���> ga?jW?o߈>��A?��
?�9O?��?�V}??��>y�N?���>�E9?+�R?[�
?͌�>'�+?�w_?�B�>}�R?bN?�8?���>��(?��?f��>^��>���>i��>�n�>�*?Ov�>�R?F�?�@?��>0˷>�M�>�_i?ޗ?X��>�/?�Ԙ>r  �r  Rr  K Kz�r  K�r  �h)Rr  tr  Rr  h�h*(h+B  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
LongStorage
qX   94889222350240qX   cpuqKNtqQ.�]q X   94889222350240qa.       �       r  �r  Rr  K ))�h)Rr  tr   Rr!  uhh)Rr"  hh)Rr#  hh)Rr$  hh)Rr%  hh)Rr&  hh)Rr'  hJ�h�hVh�G>�����h�h�G?�������h��h��ubX   4r(  h�X   5r)  hYX   6r*  h�X   7r+  h�X   8r,  h�X   9r-  hYX   10r.  h�X   11r/  h�X   12r0  h�X   13r1  hYX   14r2  h�X   15r3  h�X   16r4  h�X   17r5  hYX   18r6  h�X   19r7  h�X   20r8  h�X   21r9  hYX   22r:  h�X   23r;  h�X   24r<  h�X   25r=  hYX   26r>  h�X   27r?  h�X   28r@  h�X   29rA  hYX   30rB  h�X   31rC  h�uhJ�ubX   fc_outrD  csrc.surrogate.models.modules.fx
RegressionOutput
rE  )�rF  }rG  (hhhh)RrH  h	h)RrI  hh)RrJ  hh)RrK  hh)RrL  hh)RrM  hh)RrN  hh)RrO  X   blockrP  h)�rQ  }rR  (hhhh)RrS  h	h)RrT  hh)RrU  hh)RrV  hh)RrW  hh)RrX  hh)RrY  hh)RrZ  X   0r[  h$)�r\  }r]  (hhhh)Rr^  (h(h)h*(h+B�  ��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222249072qX   cpuqKzNtqQ.�]q X   94889222249072qa.z       T5� �ѻ��=!w�<(d�A�P�e��<1���"�퍌��V�<�l=ޕ����t�=�Žk:=s��=9�=&[�<@���>#=ҫN=�1����G%4=ţż�=uΙ�p�p��Ӿ�nd�C�G����::�=5=Ht <�@=���+m;�S�=�H��n
<bv�<�O����z�����X�ܼk� ����=��<�^=��t��=��H<Q�B�.<!ݸ<�=��ȼ�'g= B=Fg�=�^=~� ��W���廖l�<���<���Mh=�����T(<u�2��e�=��<��ϻ���<f?��%}Q=Ɓ����=���=���������<�\����;)J�]�>�-F<�O{<B����`=��=���=�9�=^й��}��)r���t���4=��=O�=[��PЁ=�bϻm5��9A;
-=SԻ�1@= �/=VEg�~�?�F��Lc*���*��������<,	-�r_  �r`  Rra  K KKz�rb  KzK�rc  �h)Rrd  tre  Rrf  �h)Rrg  �rh  Rri  h7h)h*(h+C���
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�(X   storageq ctorch
FloatStorage
qX   94889222249600qX   cpuqKNtqQ.�]q X   94889222249600qa.       *>rj  �rk  Rrl  K K�rm  K�rn  �h)Rro  trp  Rrq  �h)Rrr  �rs  Rrt  uh	h)Rru  hh)Rrv  hh)Rrw  hh)Rrx  hh)Rry  hh)Rrz  hh)Rr{  hJ�hKhVhLKubshJ�ubshJ�ubuhJ�ub.