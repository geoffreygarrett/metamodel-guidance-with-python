�csklearn.svm.classes
SVR
q )�q}q(X   kernelqX   rbfqX   degreeqKX   gammaqcnumpy.core.multiarray
scalar
qcnumpy
dtype
qX   f8q	K K�q
Rq(KX   <qNNNJ����J����K tqbC���[�q@q�qRqX   coef0qG        X   tolqG?PbM���X   CqhhC+�>5[�@q�qRqX   nuqG        X   epsilonqhhC��}�?q�qRqX	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqNX   verboseq �X   max_iterq!J����X   random_stateq"NX   _sparseq#�X   class_weight_q$cjoblib.numpy_pickle
NumpyArrayWrapper
q%)�q&}q'(X   subclassq(cnumpy
ndarray
q)X   shapeq*K �q+X   orderq,hX   dtypeq-hX
   allow_mmapq.�ubX   _gammaq/hX   support_q0h%)�q1}q2(h(h)h*M �q3h,hh-hX   i4q4K K�q5Rq6(KhNNNJ����J����K tq7bh.�ub                            	   
                                                                   !   "   #   $   %   &   '   (   )   *   +   ,   -   .   /   0   2   3   4   5   6   7   8   9   :   ;   <   =   >   @   A   B   C   D   E   F   G   I   J   K   L   M   N   O   P   Q   R   S   T   U   V   W   X   Y   Z   [   \   ]   ^   _   `   a   b   c   d   e   f   g   h   i   j   k   l   m   n   o   p   q   r   s   t   u   v   w   x   y   z   {   |   }   ~      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                         !  #  %  &  '  (  )  *  +  ,  -  .  /  0  1  2  3  4  5  6  7  8  :  ;  <  =  >  ?  @  A  B  C  D  F  G  H  J  K  L  M  O  P  Q  S  T  U  W  Y  Z  [  \  ]  ^  _  `  a  d  e  g  h  i  j  l  m  n  o  p  q  r  s  t  u  v  w  x  y  z  {  |  }  ~  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �               	  
                                         !  "  #  $  &  '  (  )  *  +  ,  -  .  /  2  3  5  6  8  9  :  ;  <  =  >  ?  X   support_vectors_q8h%)�q9}q:(h(h)h*M K�q;h,hh-hh.�ubE>>ӒW�?E������?聶_l��? dy
���?n�ǯؓ�?�彎�!�?�Vhm���?��)���?�S4��?.�Aim��?��5 �j�?E��!�?to�e_�?���M)�?���C���?�x	r�?�w%p�?���I��?��(����? �J�7�?.��$�?@��f�?�4���g�?X��7X��?�-��*�?z�G2���?�����?^KP^���?�'��K��?G>Ѓ=�?�R����?a���?�s�.�r�?M/㈏��?�>Ch���?�>�E�?ʈ }���?��M�6�?�wF9��?ؙ����?%�t߬��?��Z���?ȡ$~�F�?�-�$��?�|ߴ�?��.��?���^~�?�YIyX �?;��3G��?r�Q�he�?��!��m�?AmI�Z�?lrq%���? x/]J��?}2�//��?�9�)6�?�����?��6�j�?���u��?5X<��͑?�r	�?��e�A2�?�t8�r��?1���)�?	��i�?�6(���?2�E*	k�?��	�|W�?VYZӵ��?�	�D�?�،E�?c����?@�����?���d�?����{�?�P�B�L�?й����?|a/˳��?z4����?+/[3���?zr6���?Mn��k�?��%�?�'N2�?⽗�e��?�.W��?)H�9Ð�?鴠�J�?\�.��?���Q���?�bP\Y��?m��,�?���	�?�u(�4�?��.��?\א����?�v��3�?6�{��	�?��� i�?N����y�?����?�?K�e��?@WF^q�?p�ۙ��?�+}@��?���\��?m�Gd���?��0���?H��}<�?��o���?�4�v
�?T�����?}��(���?`��Y�?T�]��?$�dG0��?1�L�U�?x�ٚ@�?ߧm�v�?˥��j&�?ˏ��`W�?y�����?�o]����?IH�]�?K�,����?v�"G���?N�9늚�?|�(��?�#���>�?H�����?��M���?Df��?�5�1��?:�a ��?	 n��?��ǯ��?������?�ӟF���?DDm"���?M|s+Sn�?���=�?��8֦�?�����e�?��	.�?P�Ѣ�$�?�ȵ?�.�?�ZZ�;��?E+�D�K�?�j ��?,�׎[�?��m�\�?�����?&�h���?v��գ7�?l�tT���?�`��r��?����?4\S��?~���S�?x��_��?��)�u��?����?� מ��?��ٶa�?@np�<�?�2�7_,�?�iiH� �?}��{^��?35�����?e99��?� �S+��?J{��E��?
p;R�?`��n��?���\g6�?k.�˞��?W4��?v�q�9�?����?�B���0�?��
�G��?��}��?c�#���?��A���?�W�_�?�3���?X�����?h]l���?������?�l��;L�?:_y��&�?P��P,�?)�@N�2�?]{�X��?�7i�`�?{`��?F��K0��?��+p,�?�o��=�?4w�Lk�?�]��~�?R2��Z��?��T�Z�?T��;�?C镔�R�?B�3�?@������?�!�ce�?��T��?�*"�P��?�����J�?cXӁ1��?���^�?+���?�? ���s?v��~��?�mpk
�?E��HG`�?$��)v�?5�_;/f�?�pk�?H�� n�?>���t��?r���_��?=���l��?���ЖP�?D��"�?[Ɗ���?����?�)�84�?�d߱@��?e�vvg�?��4b.�?��;�5�?�"��=n�?��=Sc��?9;�@W �?�Ԓ�K�?r���	�?�rRz"�?���b	�?W,����?C<gQ���?!71��?�P�Z�u�?��⮷��?��\*�\�?C�"3�?�N��NX�?��>�2��?D/���?�t�9���?o���|�?�Cځ6��?���p6��?˥���?��l���?x�<��?<=��f`�?q7}����?ۿ,����?h�
��?{��B��?Q3:p��?ե�Q֌�? �99��?�*�e̢�?�c����?�Y��?SE�B@��?�k�|2��?
���?��H�?�?�m����?M��&c>�?���s��?M�Wϫ�?�� )3�?r�9���?Jg��\��?��fϦ�?�L��KY�?�����?����`+�?����l�?���QK��?,D�r���?d.��m�?펁���?�Q�v��?:��I	��?X߲x��?ڒ�]�{�?ª���|�?���No�?�V�����?� Qd*�?���^�(�?f)�uH��?��a��?Y���)�?"}�9���?�(U=��?M��ڰ�?W[����?��I�IJ�?�M��/�?*����?J����?�%��z�?ꠊ����?
��蘤�?�}U_��?���'��?X��*��?�!��R��?%?1��?%_S<���?��	��?ߩ��p��?A�����?��~����?HP�h�*�?���"��?����tR�?�q}�#�?н��¢?hKT���?c���Ӳ�?��]�߳�?�1m�Ԥ�?Ֆ��?�߽l��?� 0d��?����)�?8?�ι�?��$����?�]���1�?�J��K��?	Uz��?�ʶ�]�?E��N��?T�����?��{�1�?�b)��s�?�d�N^��?�4�\��?��/�a��?Z3>Z��?[58@��?�����?uv:���?�O�;�?��#�N��?��'E���?�|�.��?
���z�?�úϟ�?ܕ�����? ��P��?�G�4���?�Ix|�?�y�~Q�?���M��?
�;����?��&�]�?��C4���?=�syX�?{X%�GF�?���)I�?_��`��?3o �k�?��TH(�?|��i7�?6#^'�??����?Uu'�j�?�����?�X�Dа�?�jE���?)�!����?X[�H���?^�`u��?�����?=�:�\��?�,MK�?�ߌ"o��?kڂ|�?.�̢��?�M�h���?a��}�A�?��Dw��?���!��?k�E�?��#��?P��/���?n����X�?`Ea�d?���M��?遖:��?�A6��B�?J.���?Z�����?��8 ��?!a���?�!$%��?��{^��?�@���?4�����?���S�=�?�.�	��?F�h1U�?��k���?�����?G���?��|�?z8�	�?�Y��n�?xzݡa��?L}�}{��?�6���?Q��QQ�?"3��5��?�4&��V�?���r��?T��f2A�?|̱�ݖ�?�|�/�?F��[��?�qM��?�&�f�*�?�����J�?{��ޔ!�?ڏiy�?9�3^�k�?Βj���?K�o����?�Qs���?�^� s�?���H��?���Y�?�5 xgq?l��ѭ�?ʡ�c��?��j�d�?;d!�o�?!%�"Ʒ�?��d*��?]+t�$��?��C�ez�?��R��#�?�C��H3�?.J��r�?�ۆ��?Q
T�#3�?O>��?��|�?r,q��?�����?�7b����?�F?���?���Zt�?�p����?��Pr�;�?��g��F�?��Jh.p?_c��2�?,�1!���?o�w
B�?i�����?J���y�?'W/���?g���^'�?�;�?y7.����?�{i�l�?r�fc�?Q��!�?Y+�"��?���b�?�׀k��?0Kti8��?�x� �?i(��mf�?�����?j^FM �?�9sq���?������?D�m�R}�?6��7���?�w�Խ�?�Wt�E�?lN�9(�?�0���<�?�(���J�?D2��d%�?l��,��?���H���?N��~�?TE�t0�?��L���?f��Eg�?]Zy��o�?�cK����?��_
��?�,a�am�?�-��(Զ?�$[�N��?\WM��I�?ԭˆ6�?W����b�?�7���?$���?t�/E���?��T%u�?�$��?�!(���?�dk��?6�8#_�?�@)F=��?`�/=	��?���2�(�?U/ʷ�3�?�`@o���?ң�S��?Eʽ�^��?�EDc��? ���?�?]�%M�?P�uП��?����?N��7&�?cH� `�?��>�u5�?��e@��?4-0��?��@I�?��U;�c�?
svM��?PvK�U�?�r$Z��?P�3uAf�?��ą��?HN�����?Vw椏�?��f��w�?��T�T�?n��&���?ʼ�'��?��\�M�?+�ܶ��?���s�?�"�3���?��g6z��?7<K�C�?��a��?�j�s�@�? <�ώ��?b]Lr�?_}�O�?�SŞ֦?bYx�0�?���;��?�@�{���?�?��E�?6�[2�?���ʩ�?Q���o�?1�H�R��?�Y�g���?�� 7�S�?Q����?Tu��_G�?;8՚�?�G=-���?�5�QF��? =��N0�?Υ*���?�ur���x?Z��l)��?��d��Q�?��8f�%�?lu��?�������?��SF�T�?��6�?�p�z5�?*h���?��U����?�1���?��E6�??푵��?֌�D��?�Hۓ.��?��.zס?�Pv��?�� �Q��?J��rF�?RID���?�<Р5�?�ܭ���?�/uW��?kA\�z�?{BK'Z�?O�a��?���I�?I��� �?nB&��W�?�U'�̛�?m�%�?\�h]1��?8�׸���?�x��n��?�ׇf��?�2�'�?��;����?Yg�g���?W�?s�y�?��o5<6�?u��B�U�?.T��c�?��D	?6�?��<�?�,y�C�?1��JU��?r�JA1�?����?��5���?��Dgu�?(�ҼZ(�?0�.���?'�Jw��?���Ũ?��T��7�?����?�U��C�?��B�j�?<5[��?m�]�?3��^0M�?�&/�?e*"!���?�m1w���?6�0p�]�?�SO��?��ڑv�?��ߐ��?��*�?ֆu��?6:>P���?N߲��k�?����I��?~��Bl�?�m�x��?Oz~����?��4�#]�?��>�&4�?KIOMV��?6<�9���?�yf-t��?�Xj����?	���?qf��?�	�l���?��>����?~����n�?q���9�?v�x��C�?NP�'��?��u-���?�������?��J a�?|3����?�M{�g�?ſo���?�&��?A���L3�?���.̠�?^V��r��?7��B��?v�3����?�2�fX�?��Ř��?�b�~rT�?����R��?9�K�?\ߣ���?���9�e�?�4���5�?p��~I�?_6z����?ݥ���?�s�k!�?i-���?���)��?�f ��M�?3�Ƒ^�?�����M�?�d�i��?����?gE{4�?���p�u�?_�=���?��5���?Y��|zX�?2���{I�?t1�'�?��1���?T�!�m@�?[��^��?��"���?���t�?�H��X�?��!���?�q�+�?L���	�?f�v%�X�?`�t�?��$%"�?��  O��?Xoa8u��?�Y�S��?����*�?���Ru�?��Bl�/�?I��r��?@!*1�b�?V|֫ғ�?�h▪��?l+t1���?�v���?+���]�?v���F�?X
e�N�?۫�8��?��n��?�;�!!�?�D���I�?h�R�6�?DX��_q�?�L���?���r���?5 ��u��?.��-��?+��JD�?��vT���?2��/9K�?b�����?��1�!��?;vf����?���0ԙ�?Y`{�m�?f ����?,����?������?�mp�D��?�"�S���?P��
�&�?Oҫ�|�?|���7�?�бf�k�?R�����?$,r����?�EU�+f�?6��)��?��h�*�s?��T)]�?�"�`�&�?�4Tp��?�����?��8�;7�?���.���?�_L�N�?če���?Ҵ�deё?X�k�M�?�i1[m�?���Ѿ!�? �9bO��?2ޔ/�C�?Iڏ����?��t4,�?n70U���?a4���?SY��0�?���$��?�����?�^���N�?�?ʞϨ?&�/�8~�?������?X��ҸP�?]N�p��?;I���<�?<i����?l�i���?z���Α?AW���?ω��?��?k�#'(g�?��L�?��g@�?�i@��W�?������?�h�Z��?�.N�y��?Ӟ��5�?FQ����?W�*�`�?��YEaa�?-��qr��?�k�Y��?������?)�9��?��Ʉ2��?s�@e~�?-a%)��?�:0���?�D��#�?�w�q���?�#��\��?����Ҧ�?Ms�k�?Po�	�?�s�ݯZ�?t�����?�LJ�3�?�7s�v-w?�ߟݐ��?��n���?�YN0��?Sb�����?��I��?҉i�z�v?��aM��?�l���?�Ӝ�WH�?8c@G�H�?$�Z~"�?qFH5z?Lx�@V�?k�0Y|j�?�;^U���?R�Ij���?��7V��? ��w���?O �L��?ɨ��E{�?�ϷTَ?^��B���?B�� ��?n�����?�n3�� �?ț��;�?�9����?:C�(X��?^�6�'!�?���'�J�?�{�a���??_^q�y?�SqO�#�?�h���?�^�Y�u�?g����?루X��?r�tg�?N�e��8�?��G�&x?��Zr��?����C�?Y���B�?K�y���?@|�<�W�?���IMpy?A��b���?Ϭ�#|�w?|�$q���?�	�a���?�����?��}��?����?�K p�?|啒��?�G���x�?�m��5}�?{��[�?B�u����?¿����?w�/����?��ӛ�?{��f��?Bj�ӯQ�?t�ԓ�Z�?���pK��?Ə��W�?�LB�O\�?촘�7�?�����?�Q=Q��?�h7��?L����?^|3:h�?����[�?I1�w���?a��I���?PF2���?���|��?Ni[�?o���(_�?y�"/��?�"�CJ�?�=����?�n�|��?L�q��?K����?�q实�?^��\�6�?+�k��I�?���50�?��>���?�-�'��?N1�~�?˧�DQ+�?��3h�?������?��^p�+�?LJ+6WL�?"�L}4��?���W��?B���L�?�X�r���?�L(�S�?E�90J�?q�-Qӝ�?�R^�L�?v�;���?���E��?�u�4]�?�	�6(`�?q/%Y�?���`�?�������?������?��$����?	Jo��6�?	����C�??=t3C@�? ���C�?.�P|�?h.�@��?��Z#=>�? ��Ց}�?ۀ�`t��?F��en�?��'�j;�?��eQq��?�kj�=b�?���x�C�?>����?�hRb?�?@����?�M����?��n��`�?ƥ����?Xc�@'��?c@I�C�?�"�r(�?�O�U��?�������?B��z��?m6CF�1�?��c  �?�X�r0@�?>�U'>��?0>���?MQ�ފ��?�.$1E��?T��[΅�?�`%q���?����C�?l/�ߚ�?H���ʊ�?���3�?�-�Z�?n��-�?oА�i�?���o�?�]�֪��?��&�m�?R~�$k �?Ww��U��?���|-�?��D�?t�Zu!�?�}7p�)�?h�dGX�?�Y�}�?ђi	;n?UrX��-�?L}��c��?�腐��?K
�0O�?��P�G��?D0�t?�������?jK
�]�?t>�8�?ݢ/��C�?U�GM���?w�ź#�?�)Kϲ��?l��C�?W����2�?Iزo�Z�?���0��?����C�?G�4o��?e���zB�?�QM�c��?K.��{�?�O�샙�?\�Oe�?�w`�f��?7BT���?X
   n_support_q<h%)�q=}q>(h(h)h*K�q?h,hh-h6h.�ub        X
   dual_coef_q@h%)�qA}qB(h(h)h*KM �qCh,hh-hh.�ub��:M��S(�	6@�Q��:@�l	�v ���x^ �@��{�n��`�-J�܍J��=�A��,7#@�kq��W@m��R$@J%1w���?㕰�
�E����DB�t�]�,@�	�h�$@�M�n@(J�*T�@�gF=��+A��`�;��h^��@�"��3�c@>�@t�@�i�e��A:��"��?�$k�X@�[T5�����q'1@�8��_E@Y�N�06@\���!A@��S��64@�$����@p�<*Y*@����+@<]��@��\�A�l0�(�T"�Չy��0���
?�
 ��>�6��5&f@�ho��7@�k��	�qA�Jˡ�a^bw�	@�K~K'~�_͔�)��D���p ��Ԥ��Q@��F�|'@�c�h~>&@ϰ�t�k󿄱V�Q/��["5�4@��|1��1@��Z�@�M�� |;@�j�X��N�B�B(2@�8�l�"@��*�7(n���"����@�T��?�?���zH��?�<�qtnG�+g��Q�.�����|P���{���@4����%@��C@b�FKc@An,8�r)�3��M>0��/0�n$@�NPF3��9$���6@��z���-��e\a+@���'	@C9�VA�@ի�뻼$@T����&@Ӡ��%=�_D2�R4��#`ӛ�G��?�-@�g��7��$�3�C1��qq�!�)���:�{�Y�9���¸TQc&���¤�@ѐ���9@1��^,��?F^���c2�R��;�pE@���_�%��	�1��a���b�;��+O�jG@Kw���`�*�����7�D��)�>���4;[��b�j� @��i�_�@�3���@���qݭ!��=�m(�G�'�rfK@��9���@@F>m�����EQn��?A6�g L����p��<@�$Ǔ@%��P>�"@�zVKqmB@;	�t��#�'�ѓH�K�V����9����w�:@����0@�����Is����#@3by�R�+@l0��$�����n @�FH�*@�%s�/4��ǽӯ+@���}�@��D�U4>@o4�WgJ���r�� �����V5ۿv�D^-�A�2G,�r�)@*�G�@e�B�g�3@�����o7@����!@�v�qw�#@�7]�����*v,�p��0��Mf�^L4@�z����D�
�=z[O4�a�6PQ@M�����A@��K_���4>xZ�5��gQ��#�������@#�q����?���bF�@g���O����l| $@�����&@y0��5Q���'������'��@��PS-b-�eU�L��z�-�j"@����,@*��%���ؗ4�I$����8�H@؉�{�?G��/�� @�EnE�/Di�w�@0�+PL�"������� �Lc�W��&@���#�B��w�!Ig1@K ��(@�����@6໰�B ��z�S��A��c�Zn�񿗣�\V�½�^�q��}z�#(!�7�v��)@V�(��4�S�]b��|���i(�s��i��)@�W����?�:Q�����N�J@@�c�-v=G@v�H?(,@�/^>�5@AF���x!@G���*��VA,@�&�
�9@Y�p��C@�$u1,@8{S@	��?m���~(���3��#@r�ׅ�L�2�'LW@��dF��2@��+�8)\���*,�$@R����!@|���I4!@<cz�#@�u#�(�,����4����"u@��	:�z����+@�X[|H|%@#6D$YWG�<���,���{B�+M@�U�Cp*�?��p|�<@s�;]t�*���I��O@�6o���-���B��b@��{T��B�<Ԝ"�F�Wu�n�.�+�?�v��A��tǯ;dEſC��K��7@-�ִXe-@'�a6����!a 5@��z;u�3@\���ID@ݦ�H�h@���F�lÿP��L0�X�ה�5�n@M7��H5���Ⱦ �!@��I�L1��b�@b�1@��|�<���4D1�7@����V0@V��t`Q@7 ф{8@y��V+�%@c��D��.�7���=@�)�u��H@�L<�P�]@��4�9��J��i��s01�-@ѳ����%�����I���'�bF@
�Y8:����iF�9�Ƕ�#�U ҮIX@��Tm�@h���_�.��#T�D�2����vL;E@Gϒft�F@&�ɨ�a@��N <�9�mA�M@�����D��D�`m:/@ح�r�?�R�0U��P�r+�Ql6@�H���N���)�B��y���sX@�ї�>@ �oRfJA@��]���2@�2I"y�@�0�4��rh�2����b�W+@�_4�P2@�atƉ@�2��Ƴ�H���[*@�"��7�5@̓}��J@o���(d���(o(�26<ԗD����.TF@��\q��5��K�<m@�T�3v�c�?�|?Q��޿Q$�/Y�M��%Zt1���*+����^��X'��7|�!@�ak�"@�Q8t+]@:���P��ӵ�<@���Z�i&�A	�����0��%�N����K@��R3��!@,��&�7@u�*m�!@J���ܢ@c�ݏ�c1@�ٱ?�@��].UUC@�T��
�X�ϺG�%�'@a��޸�3��R �3i����q�4@��F�4��?�*J3@+��f@B��wt��@`�_V�*��IX���? ��ս1�"�-%��2��M��N
2����g5��b�Z*�?��;�>���}�v�?�]� å�<	��%�0a�[m�A�p�ͥ'�97��<9��gu��5����%�%�ϒ�gu�&��9$5�R��6��.�:�9 ��+�����@@��&T@ϴ7ߓD@@�~��#��K��~�0@i2 ���7��Vt@9#$@O�D/��g3��a�;3 4@@�D����D���-���1�b\i�8¡�G�@.���)0��q��4�'�|ڴ8@�����
@���mb�,�gϐOd���g,/�y@ey<���]&�<9@�\@sm�}�w>@�HıN8@���~y�[���_1@�2c��b�l��ĉ)@�ج�'@$���Ы)@w�Y�B�!@�RKc[2�l�w���M�O���@@����ʿ5�0U�D�7�F]!(@�)�u�B��g�$�\@c%���'@�}�($�-��@��Vk@����22@e����?-Vc�Xp,@�
9�� @��G� C���H!�`/��㽅d@��H\R8@�k�Ys1@�i���\E���2�(
�a�c�l/@�u.*�?@�T�_��2@I:�,�6�{ŨX����9�d�J��,��#@�!��r�0@��3;~0�E[o�9L@����j��?v�P��#@��b!3@/�C�;@n�v��@��Jh {6@���ƩOe@%q	�xC�+��3��@�á�C�����7s��F��?
��a�$`�GG�:@�KkC�Qa���b�ì @�W��V��T��UtC�Wu*�:k2�oՍ��G@T!�ZUC�?v��>Ls]@ӂC_�ga��܌�Zx&��)V#i(����� @�:\e0�m6߄(�)�9u��4�J@��rw�hC��-V0~�b@��������U�9@���}E������b�̆Γ׈$����@��r+��P@V���!>@Z�دB�@���K�]Q@��q �L��
uo��)�s��q*C$�R`4��+�m�Ŏq�q?�X���U4�4YPr��@\�^;@��0���S��f�<�+�c!��gd@w���h�+@�:Bw}�>@ΠQũ�.@1�D�ֱ=��r��@�_@`I�vI�I@�<�@_�*�x�(�s��s�2 ~�+@�J��tD0�R�K�u"�f�h����{tm�8%���k�%@$���@���1�"@�y�H�p��H�*�۶��� 8@�<�F�@�o]� �f���5���?�%	�.m@�_	��8����o4��U���R7��"���$�y3���vg$�
��(@v����@+���\@��@�D2�k�'b��?�}��v4@��\n_)@�o��+^@X
   intercept_qDh%)�qE}qF(h(h)h*K�qGh,hh-hh.�ub�4d�{K@X   probA_qHh%)�qI}qJ(h(h)h*K �qKh,hh-hh.�ubX   probB_qLh%)�qM}qN(h(h)h*K �qOh,hh-hh.�ubX   fit_status_qPK X
   shape_fit_qQM@K�qRX   _intercept_qSh%)�qT}qU(h(h)h*K�qVh,hh-hh.�ub�4d�{K@X   _dual_coef_qWh%)�qX}qY(h(h)h*KM �qZh,hh-hh.�ub��:M��S(�	6@�Q��:@�l	�v ���x^ �@��{�n��`�-J�܍J��=�A��,7#@�kq��W@m��R$@J%1w���?㕰�
�E����DB�t�]�,@�	�h�$@�M�n@(J�*T�@�gF=��+A��`�;��h^��@�"��3�c@>�@t�@�i�e��A:��"��?�$k�X@�[T5�����q'1@�8��_E@Y�N�06@\���!A@��S��64@�$����@p�<*Y*@����+@<]��@��\�A�l0�(�T"�Չy��0���
?�
 ��>�6��5&f@�ho��7@�k��	�qA�Jˡ�a^bw�	@�K~K'~�_͔�)��D���p ��Ԥ��Q@��F�|'@�c�h~>&@ϰ�t�k󿄱V�Q/��["5�4@��|1��1@��Z�@�M�� |;@�j�X��N�B�B(2@�8�l�"@��*�7(n���"����@�T��?�?���zH��?�<�qtnG�+g��Q�.�����|P���{���@4����%@��C@b�FKc@An,8�r)�3��M>0��/0�n$@�NPF3��9$���6@��z���-��e\a+@���'	@C9�VA�@ի�뻼$@T����&@Ӡ��%=�_D2�R4��#`ӛ�G��?�-@�g��7��$�3�C1��qq�!�)���:�{�Y�9���¸TQc&���¤�@ѐ���9@1��^,��?F^���c2�R��;�pE@���_�%��	�1��a���b�;��+O�jG@Kw���`�*�����7�D��)�>���4;[��b�j� @��i�_�@�3���@���qݭ!��=�m(�G�'�rfK@��9���@@F>m�����EQn��?A6�g L����p��<@�$Ǔ@%��P>�"@�zVKqmB@;	�t��#�'�ѓH�K�V����9����w�:@����0@�����Is����#@3by�R�+@l0��$�����n @�FH�*@�%s�/4��ǽӯ+@���}�@��D�U4>@o4�WgJ���r�� �����V5ۿv�D^-�A�2G,�r�)@*�G�@e�B�g�3@�����o7@����!@�v�qw�#@�7]�����*v,�p��0��Mf�^L4@�z����D�
�=z[O4�a�6PQ@M�����A@��K_���4>xZ�5��gQ��#�������@#�q����?���bF�@g���O����l| $@�����&@y0��5Q���'������'��@��PS-b-�eU�L��z�-�j"@����,@*��%���ؗ4�I$����8�H@؉�{�?G��/�� @�EnE�/Di�w�@0�+PL�"������� �Lc�W��&@���#�B��w�!Ig1@K ��(@�����@6໰�B ��z�S��A��c�Zn�񿗣�\V�½�^�q��}z�#(!�7�v��)@V�(��4�S�]b��|���i(�s��i��)@�W����?�:Q�����N�J@@�c�-v=G@v�H?(,@�/^>�5@AF���x!@G���*��VA,@�&�
�9@Y�p��C@�$u1,@8{S@	��?m���~(���3��#@r�ׅ�L�2�'LW@��dF��2@��+�8)\���*,�$@R����!@|���I4!@<cz�#@�u#�(�,����4����"u@��	:�z����+@�X[|H|%@#6D$YWG�<���,���{B�+M@�U�Cp*�?��p|�<@s�;]t�*���I��O@�6o���-���B��b@��{T��B�<Ԝ"�F�Wu�n�.�+�?�v��A��tǯ;dEſC��K��7@-�ִXe-@'�a6����!a 5@��z;u�3@\���ID@ݦ�H�h@���F�lÿP��L0�X�ה�5�n@M7��H5���Ⱦ �!@��I�L1��b�@b�1@��|�<���4D1�7@����V0@V��t`Q@7 ф{8@y��V+�%@c��D��.�7���=@�)�u��H@�L<�P�]@��4�9��J��i��s01�-@ѳ����%�����I���'�bF@
�Y8:����iF�9�Ƕ�#�U ҮIX@��Tm�@h���_�.��#T�D�2����vL;E@Gϒft�F@&�ɨ�a@��N <�9�mA�M@�����D��D�`m:/@ح�r�?�R�0U��P�r+�Ql6@�H���N���)�B��y���sX@�ї�>@ �oRfJA@��]���2@�2I"y�@�0�4��rh�2����b�W+@�_4�P2@�atƉ@�2��Ƴ�H���[*@�"��7�5@̓}��J@o���(d���(o(�26<ԗD����.TF@��\q��5��K�<m@�T�3v�c�?�|?Q��޿Q$�/Y�M��%Zt1���*+����^��X'��7|�!@�ak�"@�Q8t+]@:���P��ӵ�<@���Z�i&�A	�����0��%�N����K@��R3��!@,��&�7@u�*m�!@J���ܢ@c�ݏ�c1@�ٱ?�@��].UUC@�T��
�X�ϺG�%�'@a��޸�3��R �3i����q�4@��F�4��?�*J3@+��f@B��wt��@`�_V�*��IX���? ��ս1�"�-%��2��M��N
2����g5��b�Z*�?��;�>���}�v�?�]� å�<	��%�0a�[m�A�p�ͥ'�97��<9��gu��5����%�%�ϒ�gu�&��9$5�R��6��.�:�9 ��+�����@@��&T@ϴ7ߓD@@�~��#��K��~�0@i2 ���7��Vt@9#$@O�D/��g3��a�;3 4@@�D����D���-���1�b\i�8¡�G�@.���)0��q��4�'�|ڴ8@�����
@���mb�,�gϐOd���g,/�y@ey<���]&�<9@�\@sm�}�w>@�HıN8@���~y�[���_1@�2c��b�l��ĉ)@�ج�'@$���Ы)@w�Y�B�!@�RKc[2�l�w���M�O���@@����ʿ5�0U�D�7�F]!(@�)�u�B��g�$�\@c%���'@�}�($�-��@��Vk@����22@e����?-Vc�Xp,@�
9�� @��G� C���H!�`/��㽅d@��H\R8@�k�Ys1@�i���\E���2�(
�a�c�l/@�u.*�?@�T�_��2@I:�,�6�{ŨX����9�d�J��,��#@�!��r�0@��3;~0�E[o�9L@����j��?v�P��#@��b!3@/�C�;@n�v��@��Jh {6@���ƩOe@%q	�xC�+��3��@�á�C�����7s��F��?
��a�$`�GG�:@�KkC�Qa���b�ì @�W��V��T��UtC�Wu*�:k2�oՍ��G@T!�ZUC�?v��>Ls]@ӂC_�ga��܌�Zx&��)V#i(����� @�:\e0�m6߄(�)�9u��4�J@��rw�hC��-V0~�b@��������U�9@���}E������b�̆Γ׈$����@��r+��P@V���!>@Z�دB�@���K�]Q@��q �L��
uo��)�s��q*C$�R`4��+�m�Ŏq�q?�X���U4�4YPr��@\�^;@��0���S��f�<�+�c!��gd@w���h�+@�:Bw}�>@ΠQũ�.@1�D�ֱ=��r��@�_@`I�vI�I@�<�@_�*�x�(�s��s�2 ~�+@�J��tD0�R�K�u"�f�h����{tm�8%���k�%@$���@���1�"@�y�H�p��H�*�۶��� 8@�<�F�@�o]� �f���5���?�%	�.m@�_	��8����o4��U���R7��"���$�y3���vg$�
��(@v����@+���\@��@�D2�k�'b��?�}��v4@��\n_)@�o��+^@X   _sklearn_versionq[X   0.21.3q\ub.