�csklearn.svm.classes
SVR
q )�q}q(X   kernelqX   rbfqX   degreeqKX   gammaqcnumpy.core.multiarray
scalar
qcnumpy
dtype
qX   f8q	K K�q
Rq(KX   <qNNNJ����J����K tqbC��;%$�g@q�qRqX   coef0qG        X   tolqG?PbM���X   CqhhC/��*��@q�qRqX   nuqG        X   epsilonqhhC�vjR��?q�qRqX	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqNX   verboseq �X   max_iterq!J����X   random_stateq"NX   _sparseq#�X   class_weight_q$cjoblib.numpy_pickle
NumpyArrayWrapper
q%)�q&}q'(X   subclassq(cnumpy
ndarray
q)X   shapeq*K �q+X   orderq,hX   dtypeq-hX
   allow_mmapq.�ubX   _gammaq/hX   support_q0h%)�q1}q2(h(h)h*K-�q3h,hh-hX   i4q4K K�q5Rq6(KhNNNJ����J����K tq7bh.�ub                
                                                       "   #   '   (   )   ,   -   .   /   0   1   2   3   4   5   6   7   8   9   :   =   ?   X   support_vectors_q8h%)�q9}q:(h(h)h*K-K�q;h,hh-hh.�ub�6��?s*�u+�?�u����?c*p���?V�?Z�9�?���{��?X���@G�?.�B�E�?�8�jU(�?u)��Z�?_0=+��?������?�R��ɜ�?��yr%��?g{�B�?	z&�S�?�;�!��?/|kU�?����x��?�h
`�,�?(YtI5�?��D�f�?$M�Ӌ�?s/�pU?�?_��`.�?������?��d2h�?�U�l���?��8�_�?���?�`7 }��?
4�KG�?3T�C��?��rgXh�?���?�����L�?�'%�'x�?��\���?�61��?ۀ�Ys��?�Z�T��?�r�d��?b���?}��e��?����?��Á3��?hpP�X2�?���lM�?�k���\�?.jõDm�?"Ç�3�?�' ۸ �?
�cH�@�?�<� EA�?8'�d�?3,a*�]�?�tS3d��?��'��?��>/zC�?������?�����(�?�k��E��?�2b�4��?�x����?��r%��?\��H��?i�Wl�5�?&*JW\��?�ه�I��?�v<�ʵ?M|���? &�T�?�=�e��?R�����?"E ט��?c��C�?�!gٖ�?��4�}�?+t���?�o���?p���H��?}I|Ym��?��1k�?�L8�.�?S���L�?U�[���?r֋����?���z�?A~׳H��?�����?X
   n_support_q<h%)�q=}q>(h(h)h*K�q?h,hh-h6h.�ub        X
   dual_coef_q@h%)�qA}qB(h(h)h*KK-�qCh,hh-hh.�ubc�Q3����Q}/,�7¿7���u|ο��y�֍���@f����	R���?0��Ŋ��?���6e&п�iJs?�?f<�~`��?r���g�?ՠ��2¿4���g��?�}j��?<��o��?��а����4�<4I���y���㿠����eؿ*O��^���P� o2�?�A��gݿ�t�?��? ,�	���?L0�&W���r�/�p�����S��?�f��HQ����5�ſw;j�?ŵ���߿�	�Jd��?37��6�?5�^�"�?Nj�I<�?��+�ײ?�;�ߺ�?m�WHt2�J�dd�-����Fӿ%��Kb#ۿ��G���?,��͂�?��bp�ӿl���Iϧ�X
   intercept_qDh%)�qE}qF(h(h)h*K�qGh,hh-hh.�ub�9���?X   probA_qHh%)�qI}qJ(h(h)h*K �qKh,hh-hh.�ubX   probB_qLh%)�qM}qN(h(h)h*K �qOh,hh-hh.�ubX   fit_status_qPK X
   shape_fit_qQK@K�qRX   _intercept_qSh%)�qT}qU(h(h)h*K�qVh,hh-hh.�ub�9���?X   _dual_coef_qWh%)�qX}qY(h(h)h*KK-�qZh,hh-hh.�ubc�Q3����Q}/,�7¿7���u|ο��y�֍���@f����	R���?0��Ŋ��?���6e&п�iJs?�?f<�~`��?r���g�?ՠ��2¿4���g��?�}j��?<��o��?��а����4�<4I���y���㿠����eؿ*O��^���P� o2�?�A��gݿ�t�?��? ,�	���?L0�&W���r�/�p�����S��?�f��HQ����5�ſw;j�?ŵ���߿�	�Jd��?37��6�?5�^�"�?Nj�I<�?��+�ײ?�;�ߺ�?m�WHt2�J�dd�-����Fӿ%��Kb#ۿ��G���?,��͂�?��bp�ӿl���Iϧ�X   _sklearn_versionq[X   0.21.3q\ub.