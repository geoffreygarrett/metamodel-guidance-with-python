�csklearn.svm.classes
SVR
q )�q}q(X   kernelqX   linearqX   degreeqKX   gammaqcnumpy.core.multiarray
scalar
qcnumpy
dtype
qX   f8q	K K�q
Rq(KX   <qNNNJ����J����K tqbC R&5�g�@q�qRqX   coef0qG        X   tolqG?PbM���X   CqhhC��yg�{@q�qRqX   nuqG        X   epsilonqhhC�#�	��?q�qRqX	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqNX   verboseq �X   max_iterq!J����X   random_stateq"NX   _sparseq#�X   class_weight_q$cjoblib.numpy_pickle
NumpyArrayWrapper
q%)�q&}q'(X   subclassq(cnumpy
ndarray
q)X   shapeq*K �q+X   orderq,hX   dtypeq-hX
   allow_mmapq.�ubX   _gammaq/hX   support_q0h%)�q1}q2(h(h)h*K�q3h,hh-hX   i4q4K K�q5Rq6(KhNNNJ����J����K tq7bh.�ub                            	   
                                                   X   support_vectors_q8h%)�q9}q:(h(h)h*KK�q;h,hh-hh.�ub�2�R�?H ����?;�a��?br��-�?��a���?m)	�.��?�!l�H'�?�A�H��?.��7��?����X*�?q�5����?�����&�?����9��?���O��?(d^�"�?��DM���?�60|���?t��]/�?�2ї
b�?!��3S�?I׫bFo�?�	�)��?��@��?�nZ����?vʐ�#S�?X�0�#�?�������?�((���?I�%����?����?�����? ($�r�?M�I2h��?cngZmj�?b�4D��?H|A�q�?	�Ĥ��?�P����?�4m�ॾ?�ؼ��?r$�~��?;7?p���?�%���?�kI��%�?.>J���?u��<%��?bP[���?��3\� �?���4��?z�&���?�!�/�[�?�"�- ��?D��0���?JA"=A�?,��F�K�?W}}��?�K��?{����+�?�]|M��?8B��h�?��%(���?ޓD\>�?��<@o�?v��Z�0�?4�>�?;�̮��?D�i،$�?8�r t�?����R�?߾NS���?A�e2�?]��Ò��?��[4��?dm_��?�܍���?�	�����?�|{�F��?&�^�0��?�=���?��Zv�?3ۜ��d�?X
   n_support_q<h%)�q=}q>(h(h)h*K�q?h,hh-h6h.�ub        X
   dual_coef_q@h%)�qA}qB(h(h)h*KK�qCh,hh-hh.�ub��yg�{@��yg�{���yg�{@��yg�{@��yg�{���yg�{���	��f���yg�{@��yg�{@��yg�{���yg�{@��yg�{���yg�{���yg�{���yg�{���yg�{@N��!&/o@~�=��i@��yg�{@��yg�{�/�,��d@��yg�{���yg�{@��yg�{���yg�{@��yg�{@��yg�{�X
   intercept_qDh%)�qE}qF(h(h)h*K�qGh,hh-hh.�ub��4���@X   probA_qHh%)�qI}qJ(h(h)h*K �qKh,hh-hh.�ubX   probB_qLh%)�qM}qN(h(h)h*K �qOh,hh-hh.�ubX   fit_status_qPK X
   shape_fit_qQKK�qRX   _intercept_qSh%)�qT}qU(h(h)h*K�qVh,hh-hh.�ub��4���@X   _dual_coef_qWh%)�qX}qY(h(h)h*KK�qZh,hh-hh.�ub��yg�{@��yg�{���yg�{@��yg�{@��yg�{���yg�{���	��f���yg�{@��yg�{@��yg�{���yg�{@��yg�{���yg�{���yg�{���yg�{���yg�{@N��!&/o@~�=��i@��yg�{@��yg�{�/�,��d@��yg�{���yg�{@��yg�{���yg�{@��yg�{@��yg�{�X   _sklearn_versionq[X   0.21.3q\ub.