�csklearn.svm.classes
SVR
q )�q}q(X   kernelqX   rbfqX   degreeqKX   gammaqcnumpy.core.multiarray
scalar
qcnumpy
dtype
qX   f8q	K K�q
Rq(KX   <qNNNJ����J����K tqbC�c�:6�@q�qRqX   coef0qG        X   tolqG?PbM���X   CqhhC�)A���a@q�qRqX   nuqG        X   epsilonqhhCڕ:��?q�qRqX	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqNX   verboseq �X   max_iterq!J����X   random_stateq"NX   _sparseq#�X   class_weight_q$cjoblib.numpy_pickle
NumpyArrayWrapper
q%)�q&}q'(X   subclassq(cnumpy
ndarray
q)X   shapeq*K �q+X   orderq,hX   dtypeq-hX
   allow_mmapq.�ubX   _gammaq/hX   support_q0h%)�q1}q2(h(h)h*M��q3h,hh-hX   i4q4K K�q5Rq6(KhNNNJ����J����K tq7bh.�ub                            	   
                                                                      !   "   #   $   %   &   '   (   )   *   +   ,   -   /   0   1   2   3   4   5   6   7   8   9   :   ;   <   =   >   ?   @   A   B   C   D   E   F   G   H   I   J   K   L   M   O   P   Q   R   S   T   U   V   W   X   Y   Z   [   \   ]   ^   _   `   a   b   c   d   e   f   g   h   i   j   k   l   m   n   o   p   q   r   s   t   u   v   w   x   y   z   {   |   }   ~      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                    	  
                                         !  #  &  (  )  *  +  ,  -  .  /  0  2  3  4  5  6  7  8  9  :  ;  =  >  ?  @  C  D  F  G  H  J  K  L  N  O  Q  R  S  U  V  W  Y  Z  [  \  ]  ^  _  a  b  c  d  e  f  i  j  l  m  n  o  p  q  t  w  x  y  z  {  }  ~    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                                                         !  "  #  $  %  &  '  (  )  *  +  -  .  /  1  2  3  7  :  ;  <  =  ?  X   support_vectors_q8h%)�q9}q:(h(h)h*M�K�q;h,hh-hh.�ub��D�5�?����F�?�6��P�?ra�վ�?(����?ʾcmYy�?�H<}X��?n;^�U��?��(����?�2�o��?�iǈt�?��+AM��?#s����?+����?��~���?bVB}y�?<�4��?�_��Z��?���[Lp�?NgL��!�?R�l����?*p���?�bD?�A�?z���?�ӥw�:�?�����?�"-�F�??M�˒�?2!�_��?�X�����?̵�J�O�?���rƛ�?��U�8�?�����?P4�q���?벳�t��?�+e���?����m�?Oc)���?f���q��?�A0��x�?�4����?����ӱ�?3�?z��?��h��?r����e�? �K�q��?�U}�x�?U�)�?�Cd?m��?���3u�?-av�
�?9���Z��?q9����?Dc��u��?dމB�*�?'t�M�?�	p�p�?�ؑ�O��?86�k
��?x��2�I�? <���?~!��?�dS���?/nѥ��?����R�?l�K3-}�?	~�Ŧ��?j����q�?�-���?
�i���?�xD���?=yG^�j�?����c�?�`N�(	�?L��W���?�`��(d�?=�8�@o�?x���f��?�Q��O�?�=^����?pa�kY5�?��At�W�?. �wŊ�?��WB�V�?y�+L*�?��@��?���[9�?�N����?I��I�?L��$/��?4�F���?��S��?�2p���?0QB����?�zR:t>�?Y^he.��?�jS)@�?��y)��?��Fo�*�?�m�D�S�?s�bR�E�?#̢I1��?�cy�;��?s���Q�?����?�?�拸�? ���N�?�.����?R��;���?=b�{�?����'O�?1�1��V�?�uό�E�?ܗ���(�?f�#�i�?;$�Te�?>A���:�?�ۺ�OY�?ŚǖI��?���[��?�h�?5�����?M)�:WK�?�dy��?�tm�|�?T��?1��8ퟸ?�Mvl!%�?�Z��)$�?�3?:,z�?,��H��?ou Q�?�?,,��?���R���?���f�?s8W_3�?l�{���?�������?%�`�^�?C�qVM��?���c��?��M�KN�?qF���?ݢ�Ej�?��\6͚�?Qd\��j�?�짯�?��R���? ��P��?.�Kݣ�?`�d���?>����C�?z'.P���?�S�Q:��?�5���?:�,�!��?ܒ{y��?�������?�Д��?'xV����?z��9���?�v;I@�?:L��?W{ό}��?�%R�9.�?�T���?���3�k�?Y�����?c�_����?l��dg0�?�������?63�>��?8��J>*�?g����?h��`�{�? 1�/��?������?��J�H�?��p(��? hso�&�?t˻=�?@��4�[�?�Z���(�?
�kL��?w�ǰ��?h�Z���?D�\���?]ڋQ�`�?��xl��?�������?�!��by�?s6����?����yJ�?�e�����?�n �-�?m�+����?��YY�?�й�t��?{��QQ��?ɭ��`�?�:P;���?�Χ��?l����?�5�i���?F?ޕz�?9�uJ1�?
,��?��<���?�^��7�?���^�a?�� /j�?G���?�ka���?x�|܅�?p Q�?H����?s���a�?K����Х?+�m����?�&�<؈�?��%�Tg�?��	I�A�?H�D%���?M�ɕ��?����ٗ�?ǬG Z�?e���˔�?8数2�?����?��?@���^�?�ܶ.���?3~X���?�˯F�u�?	��FB�?�$`�+��?�Y��̾�?�=�R��?$�����?�!V:BN�?��Q)z��?���6���?���ɀ��?�W{�`�?0r@��{�?�tC��.�?������?�:����?ov[dN�?��eiC�?h�؀�?�,����?��-3��?��I�1�?�d�ݶ�?�o5�K�?�+��M�?�T+��?6��DX�?�7C�q�?�'��q�?���έ?2��.�?a��+X�?C���t��?�4[��?p�9����?�=G�[�?_���?�Tt]ly�?��Oe���?45�!�?r�N��?
�s0���?o�S�6�?`�F^*^�?�������?�q���9�?J��l:�?=��`�?��j1��?����ӫ�?;���?sݍ`���?�ݗq|G�?If5��?��	�e�?I���ob�?m+)B��?Qv�ir��?�^��e�?�2���?1՛�jk�?϶J��?�����?�Czs��?��l ��?m?���?$�[\ؼ�?H�
�x|�?{`�/��?�Gո���?��2>��?���[7�?H�sj�a�?A& ����?�C�K~��?-�AXؠ?t��}��?��y���?��r�r�?1�Q�M�?xj�����?a�L�/��?��u����?|O�@i
�?5�\����?�|-T��?�!����?0��c�x�?q�	�"�?�M�[��?��sڨ�?�`}���?�yc�?�-)���?8��4}�?�^RT��?�U�y��?��d���?밴����?�l@���?BO$���?{G�Ip�?q���?Դ�<��?aԂ�?wN�;W��?��;�#��?�?P��?(���/��?�@��	��?�Ս&�t�?���I��?�j9QuV�?�K��d%�?��u�ٲ?tU�y�J�?n�A��?Ynl:��?��U�$��?�#X>M�?�ט|ɢ�?�� �>��?Y��;��?C�E6��?8���k�?��C�;[�?*8�>{��?�����?+��a�?,d����?�6��z�?�������?�f/�4�?eMuΎ�?�$!~�?���&��?/I��2��?�Θ3	]�?�(8^���?!ai��Н?�/G�m�?}!�^'�?�-Pɫ�?����r�?��8��:�?��E�>�?��b���?�����?dǨwZ��?�����t�?�+Yc��?!w���?q�%5���?����޻�?%�Lt!!�?tQ \���?y��a���?v�tiU^�?DU�"���?XJ�Ö��?W�UH���?�L���?�gpG0�?�`'Y��?<
��~m�?d/cV�?���H�h�?���e�A�?�@Շ{�?�t7�t��?,E��T�?�xFb���?�K�ּ�?�9\:�?��
0v�?M%�uW�?�pbض�?�.r҅��?��uh��?ƍA���?� M��?[����?=w����?j�T��?����?�����r�?��U��	�?^O3�?!5Q%�Z�?��T��?qG?���?��EN�?��TO��?�K��g�?�\?X���?�Y�g[�?��fĽ	�?~�p��6�?�D�@�l�?�,�b��?e�e��?%tA��V�?��Ȯ�?~���0��?��'��?cF5����?�{]���?^��^v{�?Y�#�?����uq�?�X6��E�?�[��(��?�z�f���?������?)�X�A��?��B�Is�?z��@!=�?��ّ��?X-�?��}�G�?#�2�	�?�]�����?2+�A|$�?m���E��?Cc��6�?ҜIjM�?2{��H;�?C�G���?��"��i�?U[�%��?k�j=�?<6�L���?�������?��5x9��?�{�~�?��� 1l�?
X����?��\���?��E���?�A�p�?���/`��?+S�Bq��?j�� �?�l�y���?�����?>D:��?�	
8@�?�|��a��?E�UÃ�?C|��,.�?�r߫F<�? �&T���?��b�d��?��^��?z��.%��?g=rj��?�����?�Gj|�p�?#M6���?2����B�?O֬�F�?��iR!�?3���?�};9�?oy��O �?���Χ�?.|5a�?����?ƽ�Sn�?@4�f
�?ӮL�6Q�?����~R�?�(��ɇ�?�
pF�?�
��?�z��P�?��<���?�9�v��?��T����?��}�z�?*ƪ����?]:dYU��?6[�s
2�?�b�.�!�?�<t��?�l���?���B��?�ʼMQ9�?nUE!��?�I��Oa�?�M��A�?�b���?x�%� I�?L���F�?��?�\�?�rA&�=�?&��Ѯj�?��A�?l�G�3��?�o;���?U�vj���?ax\�P�?�Y��k��?:y�J��?�|�4R�?��ڌvg�?~�����? �G�C�?&1j1�d�?�?�IF|�?�h4�P�?�~rE�1�?bE�~���?���9�?1���?>R���X�?�s%GsK�?�n��N�?�%�$���?���g�?��7� ��?�������?���5t�?�7oM9�?��U��J�?)X.���?0A �>�?D+5�(��?�JH[���?�`��?�������?|!FfU�?͹,_�?��,�e�?.�K�?��I��S�?s��[�b�?N�m����?.��Ψ��?�*	��?�8�M�?�g�q}�?�]E0���?#ث�|�?��� ���?�D�w��?Q����?��3y���?�3����?��3�E�?-�J�?j�;���?K�y����?�5i���?<����?�������?�|�.�(�?������?vS�+�_�?�l�����?O���?��Wm8�?4��P"�?O*���?_͹�j��?7c�J�?��%؋{�?�b�&��?�u�1ֱ�?C�_d��?����4��?�Z8��?��9��@�?~Fo�Y��?��L1��?�3��o�?��G���?,�ӱ�#�?�$�썢�?�������?�P���?�-��r�?Ȅ�!���?�&���?������?���K֧�?z�����?�>4"ί?r��Rk��?�d�η�?������?��Mo��?ܺ ���?:�U34�?��o>��?l�=�$��?`��y���?S���7�?�QK�r�?�n)R�*�?�KQa�c�?�ҫA�b�?9��򇑾?{��|��?�4��]��?F����?8Y�M���?��;��?қ[��(�?痞��?|7�PE��?���l�/�?�g����?�F_ ϗ�?ӊ�����?�ӥ��?��2R{2�?��D�ۧ�?��~Hc�?�B���?�)o���?.I5���?^P�(���?W8�'���?���t0�?�~)�?.d��?��io�?���!�N�?в�N�b�?�(*��@�?�ɚ�k�?.s5���?\�E���?i]��%�?z���YL�?�>w����?Ć-���?��3N���?�4��Z�?�p���?�/,d��?Y{� �?�k�	��?R�h�.�?h��t+j�?�j�Mx��?���2���?� kǂ]�?OjM�^i�?�P���?`��O�?3a�sV=�?yxxY�%�?�ʖ���?/VU�?]��*���?���0�_�?Dn�{H��?��q�*�?��YC��?�印!�?5�>z�1�?-�#E���?�����?�^�id�?������?[�[NC�?ӌY�1��?1������?��g�qV�?�9�,Q�?�($Y�?�+G�R��?=!vus��?��@�H��?��Q�w�?-Y�!�Y�?��¾��?�O1h��?e Ŷq�?�[��v�?\��Z���?��I73�?��k�|�?p�f��+�?rO��+��?T��-N�?���?��?]�D!V��?�w�;���?T���q��?�y���i�?��g00�?�]Mm���?� 1�h�?���e�?�+���r�?^�����?v��C��?e�p��K�?υJᔺ�?=�U�?C!t���?�L@|���?�7�����?��RP��?څ����?RʽNv��?@��-��?���Z���?!�����?1;��|�?��<F�?�pP; )�?�����?AH6�av�?��;���?'
���a�?��yX8k�?�9���
�? �>x�o�?���+���?�����?ڲ���y?�5���\�?�үl��?_��̭�?�{���?�+���?��e	��?L�S�
��?.ɨ�Xs�?]��)���?�r�r
�?F3�����?��]��?4Z�Uh�?O�.�?}�-
H�?�л指�?]� t��?Y������?*�g6f�?�p��?��?�j]=���?'� ����?c
�K���?!��?�#8�?|���t�?'�&g�?T�f��?x�����?4�a@j��?��&��?��9�J��?�,H��??�<��?�?�y.�?�I�k�4�?Z�O,�?֠�5�r�?$�;Jn]�?�GiuM��?������?>��{��?̓�͂��?�M�D��?+�b�D/�?���!�?Fl����?�w	���?6�(��5�?����4�?3��b�?/�-�]�?��C+ا�?�1<����?�1T���?#��%���?��=��?';l_1�?ڲiD��?�̷��?�2u���?*�]��G�?v�����?m�I)[�?���<�?����?Dk���?�m�-I�?�B�G��?�$���?�pD����?�%5���?�
��?ɮRT3^�?�Ȯ��.�?C�\�rl�?��q�V_�?,��>�N�?�i^�@�?����M�?G�ag�/�?���Hq��?y��EN��?1��˅��?G�-�?����[(�?'"���H�??�'w�?~��>��?�\���?�6T��?� P0s
�?�0q���?3���+&�?��-Y��?��{�L1�?���54�?|��c|��?Xz%���?��?��?�U����?�[��M�?���+,L�?�),�:�?ŷU�ְ?J�O�1��?��~+�?�}�`c��?�
��?���T.�?�m S0��?����@�?iLI����?���tK��?~��e1W�?�{ 4�?y��#g�?�T�{+�?C=�4��?����+�?��Zb��?�b�����?ꖚ��	�?3qy�e\�?U>\p"�?ĸ�F���?cv��V�?�����3�?���W�?�h�+���?��u4C�?>��9�?(}����?
����?G�ùդ?�}6�2*�?� �(^�?D՞�\/�?����ph�?��\��5�?���O�Z�?�<�C��?�
r�?�~o�7�?���}�w�?g�ب�?j^v�?D%���7�?��_����?�QF��?��ތZ�?��Y��?A���.�?�#9����?��/���?0�-��?"�]���?S�/7X2�?���ܑm�?>��+�?��B�D�?�*%����?�&_�bG�?�4FdJ��?��z���?^�M��m�?����?��$��?�$���?��yL�:�??���-^?P��wN�?]v�%�?O�|�W�?���� (�?�%�����?��;�9��?��쟤��?�B�i|��?0果���?�d��+�?���4��?��ϱ�#�?ka�d���?��Daqˤ?C�r���?��ϕ��?��/t�9�?Qq��x�?�,^H�'�?f��;�[�?��в��?�a\�֧�?�eʣ��?O'�>��?*{;A\/�?}0D'��?<�j��?Y���?�?��?��'�?���
I�?�+l�4�?�\���?�-����?�S�&�?z��$��?��Et�B�?i����?��}a���?��H��>�?�q�N:�?��W��?�7���~�?( M=&B�?:y�s���?���x'�?Z�s�*�?[�7�7�?U�]�w�?#12�V��?���*Y�?�s�ѧ��?�����\�?Z]Y���?pa�1g�?���!��?� Ou��?��p�W��?�NrG�P�?�o;��(�?�E��,�?��v]��?��ds�W�?X����?��i��?E&)&�?4yǧ�?��Dj �?� N4q�?��LY���?&��y_[�? �O*{�?�̯%��?�����.�?Qd�D��?X
   n_support_q<h%)�q=}q>(h(h)h*K�q?h,hh-h6h.�ub        X
   dual_coef_q@h%)�qA}qB(h(h)h*KM��qCh,hh-hh.�ub ,#��@\�����@�\T@ӣN6��Y�?s��&M�e��?������P��Q�j.�����Vz1G��5@�88F����^���?ˬ�c��?iZx����?�Ot�Pκ�S� �}���
���?���������ʁ�@5��(Y
@�78��@/��[�-@y�����Ɲ��@b(!�I@\�ÿ' ��y�@��o�ݾ�?�,O���#��/8����h��o ��f,*�L@ .������ke2����kMk�?������P?�	�v��5K7_��࿾�\�1ͿL����?Ƣ�7�@?Š�	��'j~�+�@V�{	"�v,�[&@����M!�`����
@�6��z�;�7tn��0@tQ�%L�?�mbl8�ڿ��;M��	@��f7�����_.wT @���/��?���n��?-�h��7�?-?:��ɕ��MJ0����l @ŝ�\Uҿ�e;���꿻IO�@��b����=���?�kFK�@�����?U�?��@v��K��~4�!�����=�?�|�+p!�B#�;"@6��Tߴ�@��L��?{)jb����1��@@�3�D %���	������_�E��e
�W���i7���	@?���?E��
���ݰ��!@�}�n�?�\ݹ��?��2b��66��u*@��	%|����c��9��??9-��E@�r��s�(�S�h�����18L@�7�Q"�@702TB��?"�ooEe��������?mK�������A@~lD�.���y�8@Ə�����V+)2п�� ��? �a���
��~�n�@Yt��?���5�*t�)@��r���@��Pφ @ �wǸ�;�ع ���̓Z7�?,@d/���H�]�L�h��K@~�n�%@o;q�pj@T��0�P	@��H-��|d6z @�!�A�.��XE��@���J�@�,!M4�?�2iާܺ?֎do�@����
�n��k���.I1���IU1n���S��Re���#��@�
��R���A�D��?�0���k�?���h�:뿊��U`0@��cv�)����]��B���R�?*����=E�����?�
H�T@����Q��-�j\~3�:���@�1�o�6�?�pݽ@\�0�U��v+��@D�Ր���?��@F~�������:W)0 �@���M�?�w2�%@C#�������w�@{�<��H
�L|�<�ڿ���u @�Y�_#:�?%���0�6��o��J����@&H�ԆO@ęV�g�@�E#���>��v%@̜T-@��k`@���i���d���ҿ�w<��Z����a3׿pZ/�K@�_�/��
@oi������@50�G���Bs�7�@� �Ců�?d��*"@j�b�ɯ�?�'B�X�?���@�4p����?�O#d6@�?h���?_� �@���,�M�eL���sV(�@Ο �P�����H���"�A`�o��&@�;l�;T!�A�Iǁ�?��q���ѿ5���Q�1�.[��ZB@:���x�@� 4��7��j,��A@�+נ�u�@徢�^�?���,#l"�nd�|`@爍 ]S.@O���(	��C�4�@�G���� ��=�L#���{g�0@�@[s�*�?JĴ�B!@�!��gd���,<5���7�����ڰ���^���p'4@c\�)
����f\	@M���]�@j��+��@p#��Z����E�t8������?$�ܧ���@2��?�a��b��5C	�t�[!T�103�2�f֔d#@�6���@�oV�J<�d�g#�ms�Þ(�
�z�]� �X%U�^YL�Lx�����N+��?���P�51��n�n?@��
�0F@��"~4� ���N~�AH7�'�W=��
��:o�����̡�@h"���3@����ì@��gz=@��y;,�٪�.�h ��ٔ�@���-���(���Ţ�9`�||���5�������@��Z������B3!@�o-Ȋ�!@��������"A�@B�u
h<����Fq���y��K@�L��u#*�U�(�����8[eG��}E���]N�5ܢM�@ @�J����ٓ����A���!�/0N�Q��4һc�6@M�o��i@�F2�2@����!O�P�%#��@�(���
����8��$�Fs?�?Nă�v$@-��(@��^�Xv����-J��@���ǻ�0@��G<=2@���Dm'@�)�~X1���(��?�����cӿћy�7��?U6|� �@� \��*@|;1����?�F�y�@���La1�=2V'4��i˃�tp���>�0�@xW��@῿C�>n�&�D�㸌��X���P���3"�b��#@��W��9@��c:���q�t�������1�`�����@(�Ԧ�?}J��aM@��(KY&,�`O;X.�t�SKR𿭀� �G0@�I��C�2�$�N�#@���p��?�J-Y�e@��j����Ή\e����zv��?�x,�4@x7��,_@�	Y:@�t�*�4@[��+2�?[k�l���1�Fu��A�dl@�:|��?��-����?,㘬^@�VzVj@��'qѿ�rT�!!��ܻ�l��>���m@����� @�i3��	�iwB؍]@����ޘ
@�u�@
��/��ʶ̦��?��}�d"@��d� @=�`�?&mUO�@�j5F����1�6i��2.ߑ))�s-���7@�'�~��?��\�5ڊ}�����$@|�J�B�?J�3��	�p0':�DJ��g@*H��$e@)�рBIT�K�nS=@2��j�����PH�$�M��gEl@>%G�@;_U����? T� � �����s���x4�)�~�}5S��?ϗt�a��?X҇�{<@!�#������9p"@�<��y�'����s��1@�O�<O�?�_i/�@
S&�
����i
j@#��l�WV�%�X�8�@#E%3���?^��z��@��U�%@ �:d6�?/�h�? @9�9��#2@�f��<'@���z��@����(!@�
�6����V�#�E����=���i^�r%@6n/VN�@nQ��e~��d<8׿޿KH���1T@ޢ�o�� @�/��TU@C\�|��-~o�h�(@�w���"�;�A���V<"+�>���ډ@�l�6��޿�$ޜ�XZ@�M�!������uY<���y�L��zZ��?IEH��@Bи	�@F� �9�����[1�T�鐚/@��}����`�/�@iV$6bz0@���A�V"@�o�
1@�Lɞ?�Yɀ�=�@@�Py#*�z0�;@�u�O���?���R�j�����dF���|�1�@(�z*����鰴Nֿtt>2-���~�H@�#Tt��?�Tn��������-r���	�66���H	��'��
�Jj_@9�e�c�ۤ�Q������1��@}��$��?y���-��L��К"@���ٹ�n��"܌��X��O @+�S� @�c�b<@�L^D��@Oj�h@�vێ ����b=�O���ۓ���?ϤҪ@��^�1@�D���[ ��������:� N��[^�X��򿯆[P��D�3�鰗4@>%��;�@�k�`�+��{��F�E@���y�?��d��vt�uO@�x��7!@��׫Q�%R G@@s�&c��$@ 7�ʖ���UD����k%� )@���f��@	����3���`���l��*���ڂ#Y(���$<I�D��CX,@����S"�fN�C@X
   intercept_qDh%)�qE}qF(h(h)h*K�qGh,hh-hh.�ub6��\@X   probA_qHh%)�qI}qJ(h(h)h*K �qKh,hh-hh.�ubX   probB_qLh%)�qM}qN(h(h)h*K �qOh,hh-hh.�ubX   fit_status_qPK X
   shape_fit_qQM@K�qRX   _intercept_qSh%)�qT}qU(h(h)h*K�qVh,hh-hh.�ub6��\@X   _dual_coef_qWh%)�qX}qY(h(h)h*KM��qZh,hh-hh.�ub ,#��@\�����@�\T@ӣN6��Y�?s��&M�e��?������P��Q�j.�����Vz1G��5@�88F����^���?ˬ�c��?iZx����?�Ot�Pκ�S� �}���
���?���������ʁ�@5��(Y
@�78��@/��[�-@y�����Ɲ��@b(!�I@\�ÿ' ��y�@��o�ݾ�?�,O���#��/8����h��o ��f,*�L@ .������ke2����kMk�?������P?�	�v��5K7_��࿾�\�1ͿL����?Ƣ�7�@?Š�	��'j~�+�@V�{	"�v,�[&@����M!�`����
@�6��z�;�7tn��0@tQ�%L�?�mbl8�ڿ��;M��	@��f7�����_.wT @���/��?���n��?-�h��7�?-?:��ɕ��MJ0����l @ŝ�\Uҿ�e;���꿻IO�@��b����=���?�kFK�@�����?U�?��@v��K��~4�!�����=�?�|�+p!�B#�;"@6��Tߴ�@��L��?{)jb����1��@@�3�D %���	������_�E��e
�W���i7���	@?���?E��
���ݰ��!@�}�n�?�\ݹ��?��2b��66��u*@��	%|����c��9��??9-��E@�r��s�(�S�h�����18L@�7�Q"�@702TB��?"�ooEe��������?mK�������A@~lD�.���y�8@Ə�����V+)2п�� ��? �a���
��~�n�@Yt��?���5�*t�)@��r���@��Pφ @ �wǸ�;�ع ���̓Z7�?,@d/���H�]�L�h��K@~�n�%@o;q�pj@T��0�P	@��H-��|d6z @�!�A�.��XE��@���J�@�,!M4�?�2iާܺ?֎do�@����
�n��k���.I1���IU1n���S��Re���#��@�
��R���A�D��?�0���k�?���h�:뿊��U`0@��cv�)����]��B���R�?*����=E�����?�
H�T@����Q��-�j\~3�:���@�1�o�6�?�pݽ@\�0�U��v+��@D�Ր���?��@F~�������:W)0 �@���M�?�w2�%@C#�������w�@{�<��H
�L|�<�ڿ���u @�Y�_#:�?%���0�6��o��J����@&H�ԆO@ęV�g�@�E#���>��v%@̜T-@��k`@���i���d���ҿ�w<��Z����a3׿pZ/�K@�_�/��
@oi������@50�G���Bs�7�@� �Ců�?d��*"@j�b�ɯ�?�'B�X�?���@�4p����?�O#d6@�?h���?_� �@���,�M�eL���sV(�@Ο �P�����H���"�A`�o��&@�;l�;T!�A�Iǁ�?��q���ѿ5���Q�1�.[��ZB@:���x�@� 4��7��j,��A@�+נ�u�@徢�^�?���,#l"�nd�|`@爍 ]S.@O���(	��C�4�@�G���� ��=�L#���{g�0@�@[s�*�?JĴ�B!@�!��gd���,<5���7�����ڰ���^���p'4@c\�)
����f\	@M���]�@j��+��@p#��Z����E�t8������?$�ܧ���@2��?�a��b��5C	�t�[!T�103�2�f֔d#@�6���@�oV�J<�d�g#�ms�Þ(�
�z�]� �X%U�^YL�Lx�����N+��?���P�51��n�n?@��
�0F@��"~4� ���N~�AH7�'�W=��
��:o�����̡�@h"���3@����ì@��gz=@��y;,�٪�.�h ��ٔ�@���-���(���Ţ�9`�||���5�������@��Z������B3!@�o-Ȋ�!@��������"A�@B�u
h<����Fq���y��K@�L��u#*�U�(�����8[eG��}E���]N�5ܢM�@ @�J����ٓ����A���!�/0N�Q��4һc�6@M�o��i@�F2�2@����!O�P�%#��@�(���
����8��$�Fs?�?Nă�v$@-��(@��^�Xv����-J��@���ǻ�0@��G<=2@���Dm'@�)�~X1���(��?�����cӿћy�7��?U6|� �@� \��*@|;1����?�F�y�@���La1�=2V'4��i˃�tp���>�0�@xW��@῿C�>n�&�D�㸌��X���P���3"�b��#@��W��9@��c:���q�t�������1�`�����@(�Ԧ�?}J��aM@��(KY&,�`O;X.�t�SKR𿭀� �G0@�I��C�2�$�N�#@���p��?�J-Y�e@��j����Ή\e����zv��?�x,�4@x7��,_@�	Y:@�t�*�4@[��+2�?[k�l���1�Fu��A�dl@�:|��?��-����?,㘬^@�VzVj@��'qѿ�rT�!!��ܻ�l��>���m@����� @�i3��	�iwB؍]@����ޘ
@�u�@
��/��ʶ̦��?��}�d"@��d� @=�`�?&mUO�@�j5F����1�6i��2.ߑ))�s-���7@�'�~��?��\�5ڊ}�����$@|�J�B�?J�3��	�p0':�DJ��g@*H��$e@)�рBIT�K�nS=@2��j�����PH�$�M��gEl@>%G�@;_U����? T� � �����s���x4�)�~�}5S��?ϗt�a��?X҇�{<@!�#������9p"@�<��y�'����s��1@�O�<O�?�_i/�@
S&�
����i
j@#��l�WV�%�X�8�@#E%3���?^��z��@��U�%@ �:d6�?/�h�? @9�9��#2@�f��<'@���z��@����(!@�
�6����V�#�E����=���i^�r%@6n/VN�@nQ��e~��d<8׿޿KH���1T@ޢ�o�� @�/��TU@C\�|��-~o�h�(@�w���"�;�A���V<"+�>���ډ@�l�6��޿�$ޜ�XZ@�M�!������uY<���y�L��zZ��?IEH��@Bи	�@F� �9�����[1�T�鐚/@��}����`�/�@iV$6bz0@���A�V"@�o�
1@�Lɞ?�Yɀ�=�@@�Py#*�z0�;@�u�O���?���R�j�����dF���|�1�@(�z*����鰴Nֿtt>2-���~�H@�#Tt��?�Tn��������-r���	�66���H	��'��
�Jj_@9�e�c�ۤ�Q������1��@}��$��?y���-��L��К"@���ٹ�n��"܌��X��O @+�S� @�c�b<@�L^D��@Oj�h@�vێ ����b=�O���ۓ���?ϤҪ@��^�1@�D���[ ��������:� N��[^�X��򿯆[P��D�3�鰗4@>%��;�@�k�`�+��{��F�E@���y�?��d��vt�uO@�x��7!@��׫Q�%R G@@s�&c��$@ 7�ʖ���UD����k%� )@���f��@	����3���`���l��*���ڂ#Y(���$<I�D��CX,@����S"�fN�C@X   _sklearn_versionq[X   0.21.3q\ub.